// Simple tri-colour LED blink example.

// Correctly map pins for the iCE40UP5K SB_RGBA_DRV hard macro.

`define GREENPWM RGB0PWM
`define REDPWM   RGB1PWM
`define BLUEPWM  RGB2PWM

// taken (mostly) from
// https://github.com/im-tomu/fomu-workshop/blob/master/hdl/verilog/blink-expanded/blink.v

module top (
    // 48MHz Clock input
    // --------
    input clki,
    // LED outputs
    // --------
    output rgb0,
    output rgb1,
    output rgb2,
    // User touchable pins
    // --------
    // Connect 1-2 to enable blue LED
    input  user_1,
    output user_2,
    // Connect 3-4 to enable red LED
    output user_3,
    input  user_4,
    // USB Pins (which should be statically driven if not being used).
    // --------
    output usb_dp,
    output usb_dn,
    output usb_dp_pu
);

    // Assign USB pins to "0" so as to disconnect Fomu from
    // the host system.  Otherwise it would try to talk to
    // us over USB, which wouldn't work since we have no stack.
    assign usb_dp = 1'b0;
    assign usb_dn = 1'b0;
    assign usb_dp_pu = 1'b0;
    // Configure user pins so that we can detect the user connecting
    // 1-2 or 3-4 with conductive material.
    //
    // We do this by grounding user_2 and user_3, and configuring inputs
    // with pullups on user_1 and user_4.
    assign user_2 = 1'b0;
    assign user_3 = 1'b0;

    // Connect to system clock (with buffering)
    wire clk;
    SB_GB clk_gb (
        .USER_SIGNAL_TO_GLOBAL_BUFFER(clki),
        .GLOBAL_BUFFER_OUTPUT(clk)
    );

    // PyRTL module goes here:
    wire [3:0] colors;
    toplevel pyrtl_toplevel (
        .clk (clk),
        .in_1 (~user_1),
        .in_2 (~user_4),
        .red_o (colors[0]),
        .green_o (colors[1]),
        .blue_o (colors[2])
    );

    // Instantiate iCE40 LED driver hard logic, connecting up
    // counter state and LEDs.
    //
    // Note that it's possible to drive the LEDs directly,
    // however that is not current-limited and results in
    // overvolting the red LED.
    //
    // See also:
    // https://www.latticesemi.com/-/media/LatticeSemi/Documents/ApplicationNotes/IK/ICE40LEDDriverUsageGuide.ashx?document_id=50668
    SB_RGBA_DRV #(
        .CURRENT_MODE("0b1"),       // half current
        .RGB0_CURRENT("0b000011"),  // 4 mA
        .RGB1_CURRENT("0b000011"),  // 4 mA
        .RGB2_CURRENT("0b000011")   // 4 mA
    ) RGBA_DRIVER (
        .CURREN(1'b1),
        .RGBLEDEN(1'b1),
        .`REDPWM(colors[0]),      // Red
        .`GREENPWM(colors[1]),    // Green
        .`BLUEPWM(colors[2]),     // Blue
        .RGB0(rgb0),
        .RGB1(rgb1),
        .RGB2(rgb2)
    );

endmodule
// Generated automatically via PyRTL
// As one initial test of synthesis, map to FPGA with:
//   yosys -p "synth_xilinx -top toplevel" thisfile.v

module toplevel(clk, in_1, in_2, blue_o, green_o, red_o);
    input clk;
    input in_1;
    input in_2;
    output blue_o;
    output green_o;
    output red_o;

    reg[2:0] mem_0[31:0]; //tmp7900
    reg[3:0] mem_1[31:0]; //tmp7901
    reg[3:0] mem_2[31:0]; //tmp7902
    reg[2:0] my_calculator_ctrl = 3'd0;
    reg[3:0] my_calculator_in_x = 4'd0;
    reg[3:0] my_calculator_in_y = 4'd0;
    reg[3:0] my_calculator_out_z = 4'd0;
    reg[26:0] tmp0 = 27'd0;
    reg tmp5 = 1'd0;
    reg[7:0] tmp10 = 8'd0;
    reg[7:0] tmp11 = 8'd0;
    reg[7:0] tmp12 = 8'd0;
    reg[7:0] tmp13 = 8'd0;
    reg[7:0] tmp14 = 8'd0;
    reg[7:0] tmp15 = 8'd0;
    reg[7:0] tmp16 = 8'd0;
    reg[7:0] tmp17 = 8'd0;
    reg tmp18 = 1'd0;
    reg[4:0] tmp7899 = 5'd0;
    reg was_toggled = 1'd0;

    wire[7:0] _ver_out_tmp_0;
    wire[7:0] _ver_out_tmp_1;
    wire[7:0] _ver_out_tmp_2;
    wire[7:0] _ver_out_tmp_3;
    wire[7:0] _ver_out_tmp_4;
    wire[7:0] _ver_out_tmp_5;
    wire[7:0] _ver_out_tmp_6;
    wire[7:0] _ver_out_tmp_7;
    wire[7:0] _ver_out_tmp_8;
    wire[7:0] _ver_out_tmp_9;
    wire[7:0] _ver_out_tmp_10;
    wire[7:0] _ver_out_tmp_11;
    wire[7:0] _ver_out_tmp_12;
    wire[7:0] _ver_out_tmp_13;
    wire[7:0] _ver_out_tmp_14;
    wire[7:0] _ver_out_tmp_15;
    wire[7:0] _ver_out_tmp_16;
    wire[7:0] _ver_out_tmp_17;
    wire[7:0] _ver_out_tmp_18;
    wire[7:0] _ver_out_tmp_19;
    wire[7:0] _ver_out_tmp_20;
    wire[7:0] _ver_out_tmp_21;
    wire[7:0] _ver_out_tmp_22;
    wire[7:0] _ver_out_tmp_23;
    wire[7:0] _ver_out_tmp_24;
    wire[7:0] _ver_out_tmp_25;
    wire[7:0] _ver_out_tmp_26;
    wire[7:0] _ver_out_tmp_27;
    wire[7:0] _ver_out_tmp_28;
    wire[7:0] _ver_out_tmp_29;
    wire[7:0] _ver_out_tmp_30;
    wire[7:0] _ver_out_tmp_31;
    wire[7:0] _ver_out_tmp_32;
    wire[7:0] _ver_out_tmp_33;
    wire[7:0] _ver_out_tmp_34;
    wire[7:0] _ver_out_tmp_35;
    wire[7:0] _ver_out_tmp_36;
    wire[7:0] _ver_out_tmp_37;
    wire[7:0] _ver_out_tmp_38;
    wire[7:0] _ver_out_tmp_39;
    wire[7:0] _ver_out_tmp_40;
    wire[7:0] _ver_out_tmp_41;
    wire[7:0] _ver_out_tmp_42;
    wire[7:0] _ver_out_tmp_43;
    wire[7:0] _ver_out_tmp_44;
    wire[7:0] _ver_out_tmp_45;
    wire[7:0] _ver_out_tmp_46;
    wire[7:0] _ver_out_tmp_47;
    wire[7:0] _ver_out_tmp_48;
    wire[7:0] _ver_out_tmp_49;
    wire[7:0] _ver_out_tmp_50;
    wire[7:0] _ver_out_tmp_51;
    wire[7:0] _ver_out_tmp_52;
    wire[7:0] _ver_out_tmp_53;
    wire[7:0] _ver_out_tmp_54;
    wire[7:0] _ver_out_tmp_55;
    wire[7:0] _ver_out_tmp_56;
    wire[7:0] _ver_out_tmp_57;
    wire[7:0] _ver_out_tmp_58;
    wire[7:0] _ver_out_tmp_59;
    wire[7:0] _ver_out_tmp_60;
    wire[7:0] _ver_out_tmp_61;
    wire[7:0] _ver_out_tmp_62;
    wire[7:0] _ver_out_tmp_63;
    wire[7:0] _ver_out_tmp_64;
    wire[7:0] _ver_out_tmp_65;
    wire[7:0] _ver_out_tmp_66;
    wire[7:0] _ver_out_tmp_67;
    wire[7:0] _ver_out_tmp_68;
    wire[7:0] _ver_out_tmp_69;
    wire[7:0] _ver_out_tmp_70;
    wire[7:0] _ver_out_tmp_71;
    wire[7:0] _ver_out_tmp_72;
    wire[7:0] _ver_out_tmp_73;
    wire[7:0] _ver_out_tmp_74;
    wire[7:0] _ver_out_tmp_75;
    wire[7:0] _ver_out_tmp_76;
    wire[7:0] _ver_out_tmp_77;
    wire[7:0] _ver_out_tmp_78;
    wire[7:0] _ver_out_tmp_79;
    wire[7:0] _ver_out_tmp_80;
    wire[7:0] _ver_out_tmp_81;
    wire[7:0] _ver_out_tmp_82;
    wire[7:0] _ver_out_tmp_83;
    wire[7:0] _ver_out_tmp_84;
    wire[7:0] _ver_out_tmp_85;
    wire[7:0] _ver_out_tmp_86;
    wire[7:0] _ver_out_tmp_87;
    wire[7:0] _ver_out_tmp_88;
    wire[7:0] _ver_out_tmp_89;
    wire[7:0] _ver_out_tmp_90;
    wire[7:0] _ver_out_tmp_91;
    wire const_1_1;
    wire const_2_0;
    wire const_3_0;
    wire const_4_0;
    wire[2:0] const_5_4;
    wire[7:0] const_6_0;
    wire[7:0] const_7_2;
    wire[7:0] const_8_1;
    wire[7:0] const_9_0;
    wire[7:0] const_10_0;
    wire[7:0] const_11_0;
    wire[7:0] const_12_0;
    wire[7:0] const_13_1;
    wire const_14_0;
    wire[3:0] const_15_0;
    wire const_16_1;
    wire const_17_0;
    wire const_18_0;
    wire const_19_0;
    wire[3:0] const_20_15;
    wire const_21_1;
    wire const_22_0;
    wire[1:0] const_23_2;
    wire const_24_0;
    wire[1:0] const_25_3;
    wire const_26_0;
    wire const_27_0;
    wire const_28_0;
    wire const_29_0;
    wire const_30_0;
    wire const_31_0;
    wire[7:0] const_32_127;
    wire const_34_0;
    wire const_35_0;
    wire const_36_0;
    wire const_37_0;
    wire const_38_0;
    wire[7:0] const_39_127;
    wire const_41_0;
    wire const_42_0;
    wire const_43_0;
    wire const_44_0;
    wire const_45_0;
    wire[7:0] const_46_127;
    wire const_48_0;
    wire const_49_0;
    wire const_50_0;
    wire const_51_0;
    wire const_52_0;
    wire[7:0] const_53_127;
    wire[2:0] const_55_6;
    wire const_56_0;
    wire[2:0] const_57_7;
    wire const_58_0;
    wire[2:0] const_59_4;
    wire const_60_0;
    wire[2:0] const_61_5;
    wire const_62_0;
    wire const_63_0;
    wire const_64_0;
    wire const_65_0;
    wire const_66_0;
    wire const_67_0;
    wire const_68_0;
    wire[7:0] const_69_127;
    wire const_71_0;
    wire const_72_0;
    wire const_73_0;
    wire const_74_0;
    wire const_75_0;
    wire const_76_0;
    wire[7:0] const_77_127;
    wire const_79_0;
    wire const_80_0;
    wire const_81_0;
    wire const_82_0;
    wire const_83_0;
    wire const_84_0;
    wire[7:0] const_85_127;
    wire const_87_0;
    wire const_88_0;
    wire const_89_0;
    wire const_90_0;
    wire const_91_0;
    wire const_92_0;
    wire[7:0] const_93_127;
    wire[3:0] const_95_8;
    wire const_97_0;
    wire const_98_0;
    wire[6:0] const_99_127;
    wire const_100_0;
    wire const_102_0;
    wire const_103_0;
    wire[6:0] const_104_127;
    wire const_105_0;
    wire const_107_0;
    wire const_108_0;
    wire[6:0] const_109_127;
    wire const_110_0;
    wire const_112_0;
    wire const_113_0;
    wire[6:0] const_114_127;
    wire const_115_0;
    wire[1:0] const_116_2;
    wire const_117_0;
    wire const_118_0;
    wire const_119_0;
    wire[3:0] const_120_15;
    wire const_121_1;
    wire const_122_0;
    wire[1:0] const_123_2;
    wire const_124_0;
    wire[1:0] const_125_3;
    wire const_126_0;
    wire const_127_0;
    wire const_128_0;
    wire const_129_0;
    wire const_130_0;
    wire const_131_0;
    wire[7:0] const_132_127;
    wire const_134_0;
    wire const_135_0;
    wire const_136_0;
    wire const_137_0;
    wire const_138_0;
    wire[7:0] const_139_127;
    wire const_141_0;
    wire const_142_0;
    wire const_143_0;
    wire const_144_0;
    wire const_145_0;
    wire[7:0] const_146_127;
    wire const_148_0;
    wire const_149_0;
    wire const_150_0;
    wire const_151_0;
    wire const_152_0;
    wire[7:0] const_153_127;
    wire[2:0] const_155_6;
    wire const_156_0;
    wire[2:0] const_157_7;
    wire const_158_0;
    wire[2:0] const_159_4;
    wire const_160_0;
    wire[2:0] const_161_5;
    wire const_162_0;
    wire const_163_0;
    wire const_164_0;
    wire const_165_0;
    wire const_166_0;
    wire const_167_0;
    wire const_168_0;
    wire[7:0] const_169_127;
    wire const_171_0;
    wire const_172_0;
    wire const_173_0;
    wire const_174_0;
    wire const_175_0;
    wire const_176_0;
    wire[7:0] const_177_127;
    wire const_179_0;
    wire const_180_0;
    wire const_181_0;
    wire const_182_0;
    wire const_183_0;
    wire const_184_0;
    wire[7:0] const_185_127;
    wire const_187_0;
    wire const_188_0;
    wire const_189_0;
    wire const_190_0;
    wire const_191_0;
    wire const_192_0;
    wire[7:0] const_193_127;
    wire[3:0] const_195_8;
    wire const_197_0;
    wire const_198_0;
    wire[6:0] const_199_127;
    wire const_200_0;
    wire const_202_0;
    wire const_203_0;
    wire[6:0] const_204_127;
    wire const_205_0;
    wire const_207_0;
    wire const_208_0;
    wire[6:0] const_209_127;
    wire const_210_0;
    wire const_212_0;
    wire const_213_0;
    wire[6:0] const_214_127;
    wire const_215_0;
    wire[1:0] const_216_3;
    wire const_217_0;
    wire const_218_0;
    wire const_219_0;
    wire const_220_0;
    wire const_221_0;
    wire const_222_0;
    wire const_223_0;
    wire const_224_0;
    wire const_225_0;
    wire const_226_0;
    wire const_227_0;
    wire const_228_0;
    wire const_229_0;
    wire const_230_0;
    wire const_231_0;
    wire const_232_0;
    wire const_233_0;
    wire const_234_0;
    wire const_235_0;
    wire const_236_0;
    wire const_237_0;
    wire const_238_0;
    wire const_239_0;
    wire const_241_0;
    wire const_242_0;
    wire[6:0] const_243_127;
    wire const_244_0;
    wire const_246_0;
    wire const_247_0;
    wire[6:0] const_248_127;
    wire const_249_0;
    wire const_251_0;
    wire const_252_0;
    wire[6:0] const_253_127;
    wire const_254_0;
    wire const_256_0;
    wire const_257_0;
    wire[6:0] const_258_127;
    wire const_259_0;
    wire const_261_0;
    wire const_262_0;
    wire[6:0] const_263_127;
    wire const_264_0;
    wire const_266_0;
    wire const_267_0;
    wire[6:0] const_268_127;
    wire const_269_0;
    wire const_271_0;
    wire const_272_0;
    wire[6:0] const_273_127;
    wire const_274_0;
    wire const_276_0;
    wire const_277_0;
    wire[6:0] const_278_127;
    wire const_279_0;
    wire const_280_0;
    wire const_281_0;
    wire const_282_0;
    wire const_283_0;
    wire const_284_0;
    wire const_285_0;
    wire const_286_0;
    wire const_287_0;
    wire const_288_0;
    wire const_289_0;
    wire[3:0] const_290_15;
    wire const_291_0;
    wire const_292_0;
    wire const_293_0;
    wire[3:0] const_294_8;
    wire const_295_0;
    wire const_297_0;
    wire const_298_0;
    wire[6:0] const_299_127;
    wire const_300_0;
    wire const_302_0;
    wire const_303_0;
    wire[6:0] const_304_127;
    wire const_305_0;
    wire const_307_0;
    wire const_308_0;
    wire[6:0] const_309_127;
    wire const_310_0;
    wire const_312_0;
    wire const_313_0;
    wire[6:0] const_314_127;
    wire const_315_0;
    wire[3:0] const_316_1;
    wire const_317_0;
    wire const_318_0;
    wire const_319_0;
    wire const_320_0;
    wire const_321_0;
    wire const_322_0;
    wire[7:0] const_323_127;
    wire const_325_0;
    wire const_326_0;
    wire const_327_0;
    wire const_328_0;
    wire const_329_0;
    wire[7:0] const_330_127;
    wire const_332_0;
    wire const_333_0;
    wire const_334_0;
    wire const_335_0;
    wire const_336_0;
    wire[7:0] const_337_127;
    wire const_339_0;
    wire const_340_0;
    wire const_341_0;
    wire const_342_0;
    wire const_343_0;
    wire[7:0] const_344_127;
    wire[3:0] const_346_4;
    wire const_347_0;
    wire const_349_0;
    wire const_350_0;
    wire[6:0] const_351_127;
    wire const_352_0;
    wire const_353_0;
    wire const_354_0;
    wire const_355_0;
    wire const_356_0;
    wire const_357_0;
    wire const_358_0;
    wire[7:0] const_359_127;
    wire const_362_0;
    wire const_363_0;
    wire[6:0] const_364_127;
    wire const_365_0;
    wire const_366_0;
    wire const_367_0;
    wire const_368_0;
    wire const_369_0;
    wire const_370_0;
    wire const_371_0;
    wire[7:0] const_372_127;
    wire const_375_0;
    wire const_376_0;
    wire[6:0] const_377_127;
    wire const_378_0;
    wire const_379_0;
    wire const_380_0;
    wire const_381_0;
    wire const_382_0;
    wire const_383_0;
    wire const_384_0;
    wire[7:0] const_385_127;
    wire const_388_0;
    wire const_389_0;
    wire[6:0] const_390_127;
    wire const_391_0;
    wire const_392_0;
    wire const_393_0;
    wire const_394_0;
    wire const_395_0;
    wire const_396_0;
    wire const_397_0;
    wire[7:0] const_398_127;
    wire[3:0] const_400_6;
    wire const_401_0;
    wire[1:0] const_402_0;
    wire const_403_0;
    wire const_404_0;
    wire const_405_0;
    wire const_406_0;
    wire[7:0] const_407_127;
    wire[1:0] const_409_0;
    wire const_410_0;
    wire const_411_0;
    wire const_412_0;
    wire const_413_0;
    wire[7:0] const_414_127;
    wire[1:0] const_416_0;
    wire const_417_0;
    wire const_418_0;
    wire const_419_0;
    wire const_420_0;
    wire[7:0] const_421_127;
    wire[1:0] const_423_0;
    wire const_424_0;
    wire const_425_0;
    wire const_426_0;
    wire const_427_0;
    wire[7:0] const_428_127;
    wire[3:0] const_430_2;
    wire const_431_0;
    wire const_432_0;
    wire const_433_0;
    wire const_434_0;
    wire const_435_0;
    wire const_436_0;
    wire[7:0] const_437_127;
    wire const_439_0;
    wire const_440_0;
    wire const_441_0;
    wire const_442_0;
    wire const_443_0;
    wire[7:0] const_444_127;
    wire const_446_0;
    wire const_447_0;
    wire const_448_0;
    wire const_449_0;
    wire const_450_0;
    wire[7:0] const_451_127;
    wire const_453_0;
    wire const_454_0;
    wire const_455_0;
    wire const_456_0;
    wire const_457_0;
    wire[7:0] const_458_127;
    wire const_460_0;
    wire const_461_0;
    wire const_462_0;
    wire const_463_0;
    wire const_464_0;
    wire[7:0] const_465_127;
    wire const_467_0;
    wire const_468_0;
    wire const_469_0;
    wire const_470_0;
    wire const_471_0;
    wire[7:0] const_472_127;
    wire const_474_0;
    wire const_475_0;
    wire const_476_0;
    wire const_477_0;
    wire const_478_0;
    wire[7:0] const_479_127;
    wire const_481_0;
    wire const_482_0;
    wire const_483_0;
    wire const_484_0;
    wire const_485_0;
    wire[7:0] const_486_127;
    wire const_488_0;
    wire const_489_0;
    wire const_490_0;
    wire const_491_0;
    wire const_492_0;
    wire[7:0] const_493_127;
    wire const_495_0;
    wire const_496_0;
    wire const_497_0;
    wire const_498_0;
    wire const_499_0;
    wire[7:0] const_500_127;
    wire const_502_0;
    wire const_503_0;
    wire const_504_0;
    wire const_505_0;
    wire const_506_0;
    wire[7:0] const_507_127;
    wire const_509_0;
    wire const_510_0;
    wire const_511_0;
    wire const_512_0;
    wire const_513_0;
    wire[7:0] const_514_127;
    wire[3:0] const_516_5;
    wire const_517_1;
    wire const_519_0;
    wire const_520_0;
    wire[6:0] const_521_127;
    wire const_522_0;
    wire const_523_0;
    wire const_524_0;
    wire const_525_0;
    wire const_526_0;
    wire const_527_0;
    wire const_528_0;
    wire[7:0] const_529_127;
    wire const_532_0;
    wire const_533_0;
    wire[6:0] const_534_127;
    wire const_535_0;
    wire const_536_0;
    wire const_537_0;
    wire const_538_0;
    wire const_539_0;
    wire const_540_0;
    wire const_541_0;
    wire[7:0] const_542_127;
    wire const_545_0;
    wire const_546_0;
    wire[6:0] const_547_127;
    wire const_548_0;
    wire const_549_0;
    wire const_550_0;
    wire const_551_0;
    wire const_552_0;
    wire const_553_0;
    wire const_554_0;
    wire[7:0] const_555_127;
    wire const_558_0;
    wire const_559_0;
    wire[6:0] const_560_127;
    wire const_561_0;
    wire const_562_0;
    wire const_563_0;
    wire const_564_0;
    wire const_565_0;
    wire const_566_0;
    wire const_567_0;
    wire[7:0] const_568_127;
    wire[3:0] const_570_0;
    wire const_571_0;
    wire[3:0] const_572_0;
    wire const_573_0;
    wire const_574_1;
    wire const_576_0;
    wire const_577_0;
    wire[6:0] const_578_127;
    wire const_579_0;
    wire const_580_0;
    wire const_581_1;
    wire const_583_0;
    wire const_584_0;
    wire[6:0] const_585_127;
    wire const_586_0;
    wire const_587_0;
    wire const_588_1;
    wire const_590_0;
    wire const_591_0;
    wire[6:0] const_592_127;
    wire const_593_0;
    wire const_594_0;
    wire const_595_1;
    wire const_597_0;
    wire const_598_0;
    wire[6:0] const_599_127;
    wire const_600_0;
    wire const_601_0;
    wire const_602_1;
    wire const_604_0;
    wire const_605_0;
    wire[6:0] const_606_127;
    wire const_607_0;
    wire const_608_0;
    wire const_609_1;
    wire const_611_0;
    wire const_612_0;
    wire[6:0] const_613_127;
    wire const_614_0;
    wire const_615_0;
    wire const_616_1;
    wire const_618_0;
    wire const_619_0;
    wire[6:0] const_620_127;
    wire const_621_0;
    wire const_622_0;
    wire const_623_1;
    wire const_625_0;
    wire const_626_0;
    wire[6:0] const_627_127;
    wire const_628_0;
    wire const_629_0;
    wire[3:0] const_630_7;
    wire const_631_1;
    wire const_632_1;
    wire const_634_0;
    wire const_635_0;
    wire[6:0] const_636_127;
    wire const_637_0;
    wire const_638_0;
    wire const_639_1;
    wire const_641_0;
    wire const_642_0;
    wire[6:0] const_643_127;
    wire const_644_0;
    wire const_645_0;
    wire const_646_1;
    wire const_648_0;
    wire const_649_0;
    wire[6:0] const_650_127;
    wire const_651_0;
    wire const_652_0;
    wire const_653_1;
    wire const_655_0;
    wire const_656_0;
    wire[6:0] const_657_127;
    wire const_658_0;
    wire const_659_0;
    wire const_660_1;
    wire const_662_0;
    wire const_663_0;
    wire[6:0] const_664_127;
    wire const_665_0;
    wire const_666_0;
    wire const_667_1;
    wire const_669_0;
    wire const_670_0;
    wire[6:0] const_671_127;
    wire const_672_0;
    wire const_673_0;
    wire const_674_1;
    wire const_676_0;
    wire const_677_0;
    wire[6:0] const_678_127;
    wire const_679_0;
    wire const_680_0;
    wire const_681_1;
    wire const_683_0;
    wire const_684_0;
    wire[6:0] const_685_127;
    wire const_686_0;
    wire const_687_0;
    wire[3:0] const_688_3;
    wire const_689_1;
    wire const_690_0;
    wire const_691_0;
    wire const_692_0;
    wire const_693_0;
    wire const_694_0;
    wire[7:0] const_695_127;
    wire const_697_0;
    wire const_698_0;
    wire const_699_0;
    wire const_700_0;
    wire const_701_0;
    wire[7:0] const_702_127;
    wire const_704_0;
    wire const_705_0;
    wire const_706_0;
    wire const_707_0;
    wire const_708_0;
    wire[7:0] const_709_127;
    wire const_711_0;
    wire const_712_0;
    wire const_713_0;
    wire const_714_0;
    wire const_715_0;
    wire[7:0] const_716_127;
    wire[3:0] const_718_0;
    wire[3:0] const_719_0;
    wire const_720_0;
    wire const_721_0;
    wire const_722_0;
    wire const_723_0;
    wire const_724_0;
    wire const_725_0;
    wire const_726_0;
    wire const_727_0;
    wire const_728_0;
    wire const_729_0;
    wire const_730_0;
    wire const_731_0;
    wire const_732_0;
    wire const_733_0;
    wire const_734_0;
    wire const_735_0;
    wire const_736_0;
    wire const_737_0;
    wire const_738_0;
    wire const_739_0;
    wire const_740_0;
    wire const_741_0;
    wire const_742_0;
    wire const_743_1;
    wire const_744_0;
    wire const_745_1;
    wire const_746_0;
    wire[2:0] const_747_4;
    wire const_748_0;
    wire[3:0] const_749_15;
    wire const_750_1;
    wire const_751_0;
    wire const_756_0;
    wire const_757_0;
    wire const_758_0;
    wire const_759_0;
    wire[25:0] tmp1;
    wire[26:0] tmp2;
    wire[27:0] tmp3;
    wire[26:0] tmp4;
    wire tmp8;
    wire tmp32;
    wire[2:0] tmp34;
    wire tmp35;
    wire tmp36;
    wire tmp68;
    wire[2:0] tmp78;
    wire tmp79;
    wire[3:0] tmp87;
    wire tmp88;
    wire tmp89;
    wire tmp107;
    wire[2:0] tmp126;
    wire[3:0] tmp127;
    wire tmp128;
    wire[3:0] tmp130;
    wire tmp131;
    wire tmp132;
    wire[1:0] tmp133;
    wire tmp135;
    wire tmp136;
    wire[6:0] tmp137;
    wire[7:0] tmp138;
    wire[8:0] tmp155;
    wire tmp156;
    wire tmp157;
    wire tmp159;
    wire tmp162;
    wire tmp190;
    wire[7:0] tmp192;
    wire[6:0] tmp204;
    wire[7:0] tmp205;
    wire tmp211;
    wire tmp216;
    wire tmp217;
    wire[8:0] tmp222;
    wire tmp223;
    wire tmp224;
    wire tmp226;
    wire tmp229;
    wire tmp230;
    wire[8:0] tmp247;
    wire tmp248;
    wire tmp251;
    wire tmp253;
    wire tmp254;
    wire tmp255;
    wire tmp256;
    wire tmp257;
    wire[7:0] tmp258;
    wire[7:0] tmp259;
    wire tmp266;
    wire tmp281;
    wire tmp283;
    wire[8:0] tmp314;
    wire tmp320;
    wire[7:0] tmp325;
    wire[7:0] tmp326;
    wire tmp337;
    wire[7:0] tmp339;
    wire[8:0] tmp344;
    wire tmp348;
    wire tmp349;
    wire[8:0] tmp356;
    wire tmp358;
    wire tmp359;
    wire tmp363;
    wire tmp382;
    wire tmp385;
    wire tmp389;
    wire tmp391;
    wire[7:0] tmp392;
    wire tmp407;
    wire[3:0] tmp409;
    wire tmp410;
    wire tmp411;
    wire tmp422;
    wire tmp489;
    wire tmp501;
    wire[3:0] tmp517;
    wire tmp518;
    wire tmp521;
    wire tmp522;
    wire[8:0] tmp525;
    wire[9:0] tmp529;
    wire[8:0] tmp530;
    wire[7:0] tmp531;
    wire tmp537;
    wire tmp542;
    wire tmp543;
    wire[8:0] tmp548;
    wire tmp549;
    wire tmp552;
    wire tmp556;
    wire[8:0] tmp561;
    wire tmp562;
    wire tmp563;
    wire tmp564;
    wire tmp565;
    wire tmp568;
    wire tmp569;
    wire tmp570;
    wire tmp571;
    wire tmp589;
    wire tmp595;
    wire tmp596;
    wire[8:0] tmp601;
    wire tmp602;
    wire tmp605;
    wire tmp608;
    wire tmp610;
    wire tmp611;
    wire[7:0] tmp612;
    wire[7:0] tmp613;
    wire[8:0] tmp646;
    wire[8:0] tmp649;
    wire[9:0] tmp650;
    wire[8:0] tmp651;
    wire[7:0] tmp652;
    wire[8:0] tmp657;
    wire tmp661;
    wire tmp670;
    wire tmp673;
    wire tmp676;
    wire tmp677;
    wire[8:0] tmp682;
    wire tmp683;
    wire tmp684;
    wire tmp686;
    wire tmp689;
    wire tmp690;
    wire tmp691;
    wire tmp692;
    wire tmp701;
    wire tmp711;
    wire tmp713;
    wire tmp717;
    wire[8:0] tmp722;
    wire tmp723;
    wire tmp726;
    wire tmp728;
    wire tmp729;
    wire tmp731;
    wire tmp732;
    wire[7:0] tmp733;
    wire[7:0] tmp734;
    wire[8:0] tmp767;
    wire[8:0] tmp770;
    wire[9:0] tmp771;
    wire[8:0] tmp772;
    wire[7:0] tmp773;
    wire tmp798;
    wire[8:0] tmp803;
    wire tmp804;
    wire tmp805;
    wire tmp806;
    wire tmp807;
    wire tmp810;
    wire tmp811;
    wire tmp812;
    wire tmp813;
    wire[8:0] tmp830;
    wire tmp831;
    wire tmp838;
    wire[8:0] tmp843;
    wire tmp844;
    wire tmp847;
    wire tmp850;
    wire tmp852;
    wire tmp853;
    wire[7:0] tmp854;
    wire[7:0] tmp855;
    wire tmp858;
    wire[8:0] tmp888;
    wire[9:0] tmp892;
    wire[8:0] tmp893;
    wire[7:0] tmp894;
    wire tmp918;
    wire tmp919;
    wire[8:0] tmp924;
    wire tmp925;
    wire tmp926;
    wire tmp927;
    wire tmp928;
    wire tmp931;
    wire tmp933;
    wire tmp934;
    wire tmp942;
    wire[8:0] tmp951;
    wire tmp959;
    wire[8:0] tmp964;
    wire tmp965;
    wire tmp968;
    wire tmp971;
    wire tmp972;
    wire tmp973;
    wire tmp974;
    wire[7:0] tmp975;
    wire[7:0] tmp976;
    wire tmp997;
    wire tmp999;
    wire tmp1000;
    wire tmp1006;
    wire tmp1007;
    wire[7:0] tmp1015;
    wire tmp1025;
    wire tmp1030;
    wire tmp1056;
    wire[8:0] tmp1064;
    wire tmp1070;
    wire tmp1083;
    wire[8:0] tmp1089;
    wire tmp1103;
    wire tmp1104;
    wire tmp1107;
    wire[2:0] tmp1109;
    wire tmp1110;
    wire tmp1121;
    wire tmp1122;
    wire tmp1133;
    wire tmp1145;
    wire tmp1169;
    wire tmp1172;
    wire tmp1173;
    wire[3:0] tmp1175;
    wire tmp1176;
    wire tmp1177;
    wire tmp1188;
    wire tmp1204;
    wire[8:0] tmp1221;
    wire tmp1222;
    wire tmp1225;
    wire tmp1227;
    wire tmp1228;
    wire tmp1229;
    wire tmp1230;
    wire[7:0] tmp1232;
    wire[6:0] tmp1247;
    wire[7:0] tmp1248;
    wire tmp1260;
    wire[8:0] tmp1265;
    wire tmp1266;
    wire tmp1269;
    wire tmp1272;
    wire tmp1273;
    wire[8:0] tmp1290;
    wire tmp1291;
    wire tmp1294;
    wire tmp1295;
    wire tmp1296;
    wire tmp1297;
    wire tmp1298;
    wire tmp1299;
    wire tmp1300;
    wire[7:0] tmp1301;
    wire[7:0] tmp1302;
    wire[6:0] tmp1316;
    wire tmp1335;
    wire tmp1336;
    wire tmp1360;
    wire tmp1384;
    wire[7:0] tmp1386;
    wire tmp1392;
    wire tmp1395;
    wire tmp1396;
    wire tmp1420;
    wire[8:0] tmp1428;
    wire tmp1429;
    wire tmp1432;
    wire tmp1433;
    wire tmp1434;
    wire tmp1436;
    wire tmp1437;
    wire[7:0] tmp1439;
    wire[3:0] tmp1455;
    wire tmp1456;
    wire tmp1459;
    wire tmp1460;
    wire tmp1545;
    wire tmp1580;
    wire tmp1583;
    wire[3:0] tmp1585;
    wire tmp1586;
    wire tmp1587;
    wire[9:0] tmp1594;
    wire[8:0] tmp1595;
    wire[7:0] tmp1596;
    wire tmp1604;
    wire tmp1621;
    wire[8:0] tmp1626;
    wire tmp1627;
    wire tmp1630;
    wire tmp1633;
    wire tmp1635;
    wire tmp1636;
    wire[8:0] tmp1641;
    wire tmp1645;
    wire tmp1661;
    wire[8:0] tmp1666;
    wire tmp1667;
    wire tmp1670;
    wire tmp1671;
    wire tmp1672;
    wire tmp1673;
    wire tmp1674;
    wire tmp1675;
    wire tmp1676;
    wire[7:0] tmp1677;
    wire[7:0] tmp1678;
    wire tmp1692;
    wire tmp1694;
    wire[8:0] tmp1715;
    wire[9:0] tmp1719;
    wire[8:0] tmp1720;
    wire[7:0] tmp1721;
    wire tmp1731;
    wire tmp1746;
    wire[8:0] tmp1751;
    wire tmp1752;
    wire tmp1753;
    wire tmp1754;
    wire tmp1755;
    wire tmp1758;
    wire tmp1759;
    wire tmp1760;
    wire tmp1761;
    wire[8:0] tmp1766;
    wire tmp1770;
    wire[8:0] tmp1778;
    wire tmp1779;
    wire tmp1781;
    wire tmp1783;
    wire tmp1786;
    wire[8:0] tmp1791;
    wire tmp1792;
    wire tmp1795;
    wire tmp1798;
    wire tmp1800;
    wire tmp1801;
    wire[7:0] tmp1802;
    wire[7:0] tmp1803;
    wire tmp1820;
    wire tmp1832;
    wire tmp1833;
    wire[9:0] tmp1844;
    wire[8:0] tmp1845;
    wire[7:0] tmp1846;
    wire tmp1858;
    wire tmp1870;
    wire tmp1871;
    wire[8:0] tmp1876;
    wire tmp1877;
    wire tmp1878;
    wire tmp1880;
    wire tmp1883;
    wire tmp1884;
    wire tmp1885;
    wire tmp1886;
    wire tmp1893;
    wire tmp1907;
    wire tmp1911;
    wire[8:0] tmp1916;
    wire tmp1917;
    wire tmp1920;
    wire tmp1922;
    wire tmp1923;
    wire tmp1925;
    wire tmp1926;
    wire[7:0] tmp1927;
    wire[7:0] tmp1928;
    wire tmp1953;
    wire[8:0] tmp1968;
    wire[9:0] tmp1969;
    wire[8:0] tmp1970;
    wire[7:0] tmp1971;
    wire tmp1996;
    wire[8:0] tmp2001;
    wire tmp2002;
    wire tmp2003;
    wire tmp2004;
    wire tmp2005;
    wire tmp2008;
    wire tmp2010;
    wire tmp2011;
    wire tmp2019;
    wire tmp2036;
    wire[8:0] tmp2041;
    wire tmp2042;
    wire tmp2045;
    wire tmp2048;
    wire tmp2049;
    wire tmp2050;
    wire tmp2051;
    wire[7:0] tmp2052;
    wire[7:0] tmp2053;
    wire tmp2081;
    wire tmp2088;
    wire tmp2089;
    wire tmp2111;
    wire tmp2132;
    wire tmp2167;
    wire tmp2169;
    wire tmp2195;
    wire[2:0] tmp2198;
    wire tmp2199;
    wire tmp2224;
    wire[8:0] tmp2229;
    wire tmp2230;
    wire tmp2236;
    wire tmp2249;
    wire tmp2250;
    wire tmp2258;
    wire[6:0] tmp2265;
    wire tmp2274;
    wire tmp2275;
    wire tmp2276;
    wire tmp2311;
    wire tmp2323;
    wire tmp2336;
    wire tmp2337;
    wire tmp2355;
    wire tmp2362;
    wire tmp2363;
    wire tmp2376;
    wire tmp2379;
    wire tmp2380;
    wire tmp2384;
    wire tmp2387;
    wire tmp2388;
    wire tmp2399;
    wire tmp2400;
    wire tmp2401;
    wire tmp2412;
    wire tmp2413;
    wire tmp2414;
    wire tmp2415;
    wire tmp2416;
    wire tmp2417;
    wire tmp2418;
    wire tmp2419;
    wire tmp2442;
    wire tmp2455;
    wire[8:0] tmp2481;
    wire[7:0] tmp2482;
    wire[8:0] tmp2500;
    wire[7:0] tmp2501;
    wire tmp2512;
    wire[8:0] tmp2516;
    wire[7:0] tmp2520;
    wire tmp2532;
    wire[7:0] tmp2539;
    wire tmp2549;
    wire[7:0] tmp2558;
    wire[8:0] tmp2573;
    wire[7:0] tmp2577;
    wire tmp2585;
    wire tmp2589;
    wire[8:0] tmp2595;
    wire[7:0] tmp2596;
    wire tmp2613;
    wire[8:0] tmp2624;
    wire tmp2632;
    wire tmp2633;
    wire tmp2634;
    wire tmp2659;
    wire tmp2660;
    wire tmp2671;
    wire tmp2745;
    wire tmp2748;
    wire tmp2749;
    wire tmp2753;
    wire tmp2764;
    wire tmp2787;
    wire tmp2800;
    wire tmp2801;
    wire tmp2895;
    wire[6:0] tmp2918;
    wire tmp2919;
    wire[7:0] tmp2921;
    wire[8:0] tmp2924;
    wire tmp2925;
    wire tmp2927;
    wire tmp2928;
    wire tmp2931;
    wire tmp2932;
    wire tmp2933;
    wire tmp2935;
    wire[7:0] tmp2937;
    wire[8:0] tmp2940;
    wire tmp2941;
    wire tmp2944;
    wire tmp2947;
    wire tmp2948;
    wire tmp2949;
    wire tmp2950;
    wire[8:0] tmp2957;
    wire tmp2958;
    wire tmp2959;
    wire tmp2960;
    wire tmp2961;
    wire tmp2964;
    wire tmp2965;
    wire tmp2966;
    wire tmp2967;
    wire[6:0] tmp2968;
    wire[8:0] tmp2974;
    wire tmp2975;
    wire tmp2977;
    wire tmp2978;
    wire tmp2981;
    wire tmp2982;
    wire tmp2983;
    wire tmp2984;
    wire tmp3054;
    wire[7:0] tmp3062;
    wire tmp3079;
    wire tmp3081;
    wire[7:0] tmp3083;
    wire tmp3115;
    wire tmp3150;
    wire tmp3222;
    wire[6:0] tmp3241;
    wire[8:0] tmp3259;
    wire tmp3261;
    wire tmp3279;
    wire[8:0] tmp3284;
    wire tmp3285;
    wire tmp3290;
    wire tmp3293;
    wire[7:0] tmp3316;
    wire tmp3337;
    wire tmp3364;
    wire tmp3367;
    wire tmp3368;
    wire[7:0] tmp3369;
    wire[7:0] tmp3370;
    wire tmp3387;
    wire[8:0] tmp3395;
    wire tmp3399;
    wire tmp3400;
    wire tmp3401;
    wire tmp3408;
    wire tmp3411;
    wire tmp3415;
    wire tmp3424;
    wire tmp3427;
    wire[8:0] tmp3432;
    wire tmp3436;
    wire tmp3439;
    wire[7:0] tmp3444;
    wire tmp3470;
    wire tmp3489;
    wire[8:0] tmp3494;
    wire tmp3497;
    wire tmp3512;
    wire tmp3513;
    wire tmp3514;
    wire[7:0] tmp3518;
    wire tmp3543;
    wire tmp3544;
    wire tmp3546;
    wire tmp3547;
    wire tmp3548;
    wire tmp3552;
    wire tmp3555;
    wire tmp3558;
    wire tmp3559;
    wire tmp3560;
    wire tmp3561;
    wire tmp3566;
    wire tmp3567;
    wire tmp3568;
    wire tmp3571;
    wire tmp3572;
    wire tmp3573;
    wire tmp3574;
    wire[8:0] tmp3577;
    wire tmp3581;
    wire tmp3584;
    wire tmp3585;
    wire tmp3586;
    wire tmp3587;
    wire[8:0] tmp3594;
    wire tmp3595;
    wire tmp3596;
    wire tmp3598;
    wire tmp3601;
    wire tmp3602;
    wire[8:0] tmp3609;
    wire tmp3610;
    wire tmp3611;
    wire tmp3612;
    wire tmp3613;
    wire tmp3616;
    wire tmp3617;
    wire[6:0] tmp3618;
    wire[8:0] tmp3624;
    wire tmp3625;
    wire tmp3628;
    wire tmp3631;
    wire tmp3632;
    wire[8:0] tmp3639;
    wire tmp3640;
    wire tmp3641;
    wire tmp3643;
    wire tmp3646;
    wire tmp3647;
    wire tmp3701;
    wire tmp3702;
    wire[8:0] tmp3708;
    wire[9:0] tmp3711;
    wire tmp3712;
    wire[8:0] tmp3722;
    wire tmp3728;
    wire tmp3735;
    wire tmp3740;
    wire tmp3741;
    wire tmp3742;
    wire[8:0] tmp3747;
    wire tmp3749;
    wire tmp3751;
    wire tmp3754;
    wire tmp3757;
    wire tmp3764;
    wire tmp3778;
    wire tmp3788;
    wire tmp3794;
    wire tmp3795;
    wire tmp3796;
    wire tmp3797;
    wire[7:0] tmp3799;
    wire[8:0] tmp3842;
    wire[1:0] tmp3844;
    wire tmp3846;
    wire[8:0] tmp3856;
    wire tmp3857;
    wire tmp3860;
    wire tmp3874;
    wire tmp3875;
    wire tmp3876;
    wire tmp3885;
    wire tmp3888;
    wire tmp3890;
    wire tmp3891;
    wire[9:0] tmp3908;
    wire tmp3912;
    wire tmp3913;
    wire tmp3915;
    wire tmp3916;
    wire tmp3922;
    wire tmp3925;
    wire tmp3926;
    wire tmp3927;
    wire tmp3931;
    wire[7:0] tmp3933;
    wire[8:0] tmp3976;
    wire tmp3991;
    wire tmp3994;
    wire[9:0] tmp4002;
    wire tmp4006;
    wire tmp4007;
    wire[8:0] tmp4015;
    wire tmp4016;
    wire tmp4019;
    wire tmp4022;
    wire tmp4024;
    wire tmp4025;
    wire tmp4037;
    wire[8:0] tmp4041;
    wire[9:0] tmp4042;
    wire tmp4045;
    wire tmp4046;
    wire tmp4050;
    wire tmp4056;
    wire tmp4059;
    wire tmp4061;
    wire tmp4062;
    wire tmp4063;
    wire tmp4064;
    wire tmp4065;
    wire[7:0] tmp4067;
    wire[8:0] tmp4109;
    wire[8:0] tmp4110;
    wire[9:0] tmp4116;
    wire[9:0] tmp4118;
    wire[7:0] tmp4119;
    wire tmp4125;
    wire tmp4128;
    wire[9:0] tmp4136;
    wire tmp4143;
    wire tmp4144;
    wire tmp4156;
    wire tmp4157;
    wire tmp4158;
    wire tmp4159;
    wire[9:0] tmp4176;
    wire tmp4180;
    wire tmp4183;
    wire tmp4184;
    wire[8:0] tmp4189;
    wire tmp4190;
    wire tmp4193;
    wire tmp4194;
    wire tmp4196;
    wire tmp4198;
    wire[7:0] tmp4200;
    wire[7:0] tmp4201;
    wire tmp4218;
    wire[8:0] tmp4222;
    wire tmp4223;
    wire tmp4226;
    wire tmp4229;
    wire[8:0] tmp4232;
    wire tmp4233;
    wire tmp4236;
    wire tmp4239;
    wire tmp4240;
    wire[8:0] tmp4243;
    wire tmp4244;
    wire tmp4247;
    wire tmp4250;
    wire tmp4251;
    wire[8:0] tmp4254;
    wire tmp4255;
    wire tmp4258;
    wire tmp4261;
    wire tmp4262;
    wire tmp4280;
    wire tmp4358;
    wire tmp4362;
    wire[8:0] tmp4465;
    wire tmp4466;
    wire tmp4469;
    wire tmp4472;
    wire[5:0] tmp4473;
    wire[7:0] tmp4474;
    wire tmp4483;
    wire tmp4486;
    wire[8:0] tmp4491;
    wire tmp4492;
    wire tmp4495;
    wire tmp4498;
    wire tmp4499;
    wire tmp4505;
    wire[8:0] tmp4516;
    wire tmp4517;
    wire tmp4520;
    wire tmp4521;
    wire tmp4522;
    wire tmp4523;
    wire tmp4524;
    wire tmp4525;
    wire tmp4526;
    wire[7:0] tmp4527;
    wire[7:0] tmp4528;
    wire[8:0] tmp4531;
    wire tmp4532;
    wire tmp4535;
    wire tmp4536;
    wire tmp4537;
    wire tmp4538;
    wire tmp4539;
    wire[8:0] tmp4542;
    wire tmp4546;
    wire tmp4547;
    wire tmp4549;
    wire tmp4550;
    wire[5:0] tmp4551;
    wire[7:0] tmp4552;
    wire tmp4558;
    wire tmp4561;
    wire tmp4564;
    wire[8:0] tmp4569;
    wire tmp4570;
    wire tmp4571;
    wire tmp4572;
    wire tmp4573;
    wire tmp4576;
    wire tmp4577;
    wire tmp4589;
    wire[8:0] tmp4594;
    wire tmp4595;
    wire tmp4598;
    wire tmp4601;
    wire tmp4602;
    wire tmp4603;
    wire tmp4604;
    wire[7:0] tmp4605;
    wire[7:0] tmp4606;
    wire[8:0] tmp4609;
    wire tmp4610;
    wire tmp4613;
    wire tmp4614;
    wire tmp4615;
    wire tmp4616;
    wire tmp4617;
    wire[8:0] tmp4620;
    wire tmp4621;
    wire tmp4624;
    wire tmp4627;
    wire tmp4628;
    wire[5:0] tmp4629;
    wire[7:0] tmp4630;
    wire tmp4642;
    wire[8:0] tmp4647;
    wire tmp4648;
    wire tmp4651;
    wire tmp4654;
    wire tmp4655;
    wire[8:0] tmp4660;
    wire[8:0] tmp4672;
    wire tmp4673;
    wire tmp4676;
    wire tmp4677;
    wire tmp4678;
    wire tmp4679;
    wire tmp4680;
    wire tmp4681;
    wire tmp4682;
    wire[7:0] tmp4683;
    wire[7:0] tmp4684;
    wire[8:0] tmp4687;
    wire tmp4688;
    wire tmp4691;
    wire tmp4692;
    wire tmp4693;
    wire tmp4694;
    wire tmp4695;
    wire tmp4699;
    wire tmp4702;
    wire tmp4703;
    wire tmp4705;
    wire tmp4706;
    wire[5:0] tmp4707;
    wire[7:0] tmp4708;
    wire tmp4717;
    wire[8:0] tmp4725;
    wire tmp4726;
    wire tmp4727;
    wire tmp4729;
    wire tmp4732;
    wire tmp4733;
    wire tmp4745;
    wire[8:0] tmp4750;
    wire tmp4751;
    wire tmp4754;
    wire tmp4756;
    wire tmp4757;
    wire tmp4758;
    wire tmp4759;
    wire tmp4760;
    wire[7:0] tmp4761;
    wire[7:0] tmp4762;
    wire[8:0] tmp4765;
    wire tmp4766;
    wire tmp4769;
    wire tmp4770;
    wire tmp4771;
    wire tmp4772;
    wire tmp4773;
    wire tmp4780;
    wire tmp4796;
    wire tmp4798;
    wire[6:0] tmp4848;
    wire tmp4877;
    wire tmp4931;
    wire tmp5036;
    wire tmp5077;
    wire tmp5081;
    wire[7:0] tmp5129;
    wire[8:0] tmp5134;
    wire tmp5135;
    wire tmp5150;
    wire tmp5154;
    wire tmp5175;
    wire[7:0] tmp5182;
    wire[7:0] tmp5183;
    wire[8:0] tmp5215;
    wire[8:0] tmp5227;
    wire tmp5228;
    wire tmp5229;
    wire tmp5241;
    wire tmp5244;
    wire tmp5253;
    wire tmp5256;
    wire tmp5259;
    wire[6:0] tmp5290;
    wire[7:0] tmp5291;
    wire[8:0] tmp5308;
    wire tmp5310;
    wire tmp5315;
    wire tmp5322;
    wire tmp5334;
    wire tmp5341;
    wire tmp5342;
    wire tmp5343;
    wire[7:0] tmp5372;
    wire[7:0] tmp5375;
    wire[8:0] tmp5377;
    wire tmp5384;
    wire tmp5390;
    wire tmp5391;
    wire tmp5404;
    wire tmp5406;
    wire tmp5418;
    wire tmp5424;
    wire[7:0] tmp5425;
    wire[6:0] tmp5452;
    wire[7:0] tmp5453;
    wire tmp5459;
    wire[8:0] tmp5470;
    wire tmp5471;
    wire tmp5473;
    wire tmp5474;
    wire tmp5477;
    wire tmp5478;
    wire[8:0] tmp5483;
    wire[8:0] tmp5495;
    wire tmp5496;
    wire tmp5499;
    wire tmp5500;
    wire tmp5502;
    wire tmp5503;
    wire tmp5504;
    wire tmp5505;
    wire[7:0] tmp5506;
    wire[7:0] tmp5507;
    wire[8:0] tmp5510;
    wire tmp5511;
    wire tmp5514;
    wire tmp5515;
    wire tmp5516;
    wire tmp5517;
    wire tmp5530;
    wire tmp5537;
    wire tmp5543;
    wire[8:0] tmp5549;
    wire tmp5553;
    wire tmp5568;
    wire tmp5569;
    wire tmp5571;
    wire[8:0] tmp5576;
    wire tmp5577;
    wire tmp5580;
    wire tmp5581;
    wire tmp5582;
    wire tmp5583;
    wire tmp5584;
    wire[6:0] tmp5585;
    wire[7:0] tmp5586;
    wire tmp5598;
    wire[8:0] tmp5603;
    wire tmp5604;
    wire tmp5607;
    wire tmp5610;
    wire tmp5611;
    wire tmp5620;
    wire[8:0] tmp5628;
    wire tmp5629;
    wire tmp5632;
    wire tmp5633;
    wire tmp5634;
    wire tmp5635;
    wire tmp5636;
    wire tmp5637;
    wire tmp5638;
    wire[7:0] tmp5639;
    wire[7:0] tmp5640;
    wire[8:0] tmp5643;
    wire tmp5644;
    wire tmp5647;
    wire tmp5648;
    wire tmp5649;
    wire tmp5650;
    wire tmp5651;
    wire[6:0] tmp5652;
    wire tmp5677;
    wire tmp5678;
    wire[8:0] tmp5683;
    wire tmp5685;
    wire tmp5686;
    wire[8:0] tmp5695;
    wire tmp5703;
    wire[8:0] tmp5710;
    wire tmp5711;
    wire tmp5713;
    wire tmp5714;
    wire tmp5715;
    wire tmp5716;
    wire tmp5717;
    wire tmp5718;
    wire[6:0] tmp5719;
    wire[7:0] tmp5720;
    wire[8:0] tmp5725;
    wire[8:0] tmp5737;
    wire tmp5738;
    wire tmp5741;
    wire tmp5744;
    wire tmp5745;
    wire[8:0] tmp5750;
    wire tmp5754;
    wire[8:0] tmp5762;
    wire tmp5763;
    wire tmp5766;
    wire tmp5767;
    wire tmp5768;
    wire tmp5769;
    wire tmp5770;
    wire tmp5771;
    wire tmp5772;
    wire[7:0] tmp5773;
    wire[7:0] tmp5774;
    wire[8:0] tmp5777;
    wire tmp5778;
    wire tmp5781;
    wire tmp5782;
    wire tmp5783;
    wire tmp5784;
    wire tmp5785;
    wire tmp5793;
    wire tmp5835;
    wire[7:0] tmp5840;
    wire[8:0] tmp5844;
    wire tmp5845;
    wire tmp5848;
    wire tmp5849;
    wire tmp5850;
    wire tmp5851;
    wire tmp5852;
    wire[6:0] tmp5853;
    wire[7:0] tmp5854;
    wire[8:0] tmp5859;
    wire[8:0] tmp5871;
    wire tmp5872;
    wire tmp5873;
    wire tmp5875;
    wire tmp5878;
    wire tmp5879;
    wire tmp5887;
    wire tmp5888;
    wire[8:0] tmp5896;
    wire tmp5897;
    wire tmp5900;
    wire tmp5902;
    wire tmp5903;
    wire tmp5904;
    wire tmp5905;
    wire tmp5906;
    wire[7:0] tmp5907;
    wire[7:0] tmp5908;
    wire[8:0] tmp5911;
    wire tmp5912;
    wire tmp5915;
    wire tmp5916;
    wire tmp5917;
    wire tmp5918;
    wire tmp5919;
    wire[6:0] tmp5920;
    wire[8:0] tmp5938;
    wire tmp5942;
    wire tmp5945;
    wire tmp5952;
    wire[8:0] tmp5963;
    wire tmp5964;
    wire tmp5972;
    wire[8:0] tmp5978;
    wire tmp5979;
    wire tmp5982;
    wire tmp5983;
    wire tmp5984;
    wire tmp5985;
    wire tmp5986;
    wire tmp6009;
    wire tmp6025;
    wire tmp6030;
    wire[1:0] tmp6070;
    wire[9:0] tmp6074;
    wire[10:0] tmp6075;
    wire[9:0] tmp6076;
    wire[7:0] tmp6077;
    wire tmp6086;
    wire tmp6089;
    wire[9:0] tmp6094;
    wire tmp6098;
    wire tmp6108;
    wire tmp6116;
    wire tmp6123;
    wire tmp6126;
    wire tmp6129;
    wire[9:0] tmp6134;
    wire tmp6135;
    wire tmp6140;
    wire tmp6141;
    wire tmp6142;
    wire[8:0] tmp6147;
    wire tmp6151;
    wire tmp6153;
    wire[7:0] tmp6158;
    wire tmp6209;
    wire tmp6210;
    wire[9:0] tmp6219;
    wire[9:0] tmp6222;
    wire[10:0] tmp6223;
    wire[9:0] tmp6224;
    wire[7:0] tmp6225;
    wire[9:0] tmp6242;
    wire tmp6243;
    wire tmp6246;
    wire[8:0] tmp6255;
    wire tmp6256;
    wire[8:0] tmp6270;
    wire tmp6271;
    wire tmp6277;
    wire tmp6283;
    wire[8:0] tmp6295;
    wire tmp6302;
    wire tmp6303;
    wire tmp6304;
    wire[7:0] tmp6306;
    wire tmp6327;
    wire tmp6353;
    wire tmp6356;
    wire tmp6358;
    wire[1:0] tmp6366;
    wire[9:0] tmp6367;
    wire[9:0] tmp6370;
    wire[10:0] tmp6371;
    wire[9:0] tmp6372;
    wire[7:0] tmp6373;
    wire tmp6385;
    wire[7:0] tmp6387;
    wire tmp6391;
    wire tmp6397;
    wire tmp6398;
    wire tmp6405;
    wire tmp6419;
    wire tmp6431;
    wire tmp6437;
    wire[8:0] tmp6443;
    wire[7:0] tmp6454;
    wire tmp6506;
    wire[1:0] tmp6514;
    wire[9:0] tmp6515;
    wire tmp6516;
    wire[10:0] tmp6519;
    wire tmp6533;
    wire tmp6539;
    wire tmp6542;
    wire tmp6544;
    wire[8:0] tmp6551;
    wire tmp6552;
    wire tmp6555;
    wire[8:0] tmp6566;
    wire tmp6567;
    wire tmp6573;
    wire tmp6579;
    wire tmp6597;
    wire tmp6601;
    wire tmp6653;
    wire tmp6665;
    wire tmp6680;
    wire[8:0] tmp6732;
    wire[8:0] tmp6738;
    wire tmp6740;
    wire[9:0] tmp6753;
    wire tmp6754;
    wire tmp6755;
    wire tmp6756;
    wire tmp6757;
    wire tmp6759;
    wire tmp6760;
    wire tmp6761;
    wire tmp6762;
    wire tmp6763;
    wire[8:0] tmp6771;
    wire[8:0] tmp6772;
    wire tmp6774;
    wire[9:0] tmp6787;
    wire tmp6788;
    wire tmp6789;
    wire tmp6790;
    wire tmp6791;
    wire tmp6792;
    wire tmp6794;
    wire tmp6795;
    wire tmp6798;
    wire[8:0] tmp6816;
    wire[8:0] tmp6818;
    wire[8:0] tmp6819;
    wire[9:0] tmp6822;
    wire tmp6823;
    wire tmp6824;
    wire tmp6825;
    wire tmp6826;
    wire tmp6828;
    wire tmp6829;
    wire tmp6830;
    wire tmp6832;
    wire[8:0] tmp6841;
    wire tmp6844;
    wire[8:0] tmp6848;
    wire[8:0] tmp6853;
    wire[9:0] tmp6857;
    wire tmp6858;
    wire tmp6859;
    wire tmp6860;
    wire tmp6861;
    wire tmp6862;
    wire tmp6864;
    wire tmp6865;
    wire tmp6942;
    wire tmp6951;
    wire tmp6991;
    wire tmp7009;
    wire tmp7026;
    wire tmp7027;
    wire[8:0] tmp7034;
    wire[8:0] tmp7036;
    wire[7:0] tmp7038;
    wire tmp7039;
    wire[8:0] tmp7041;
    wire[8:0] tmp7052;
    wire[8:0] tmp7053;
    wire[9:0] tmp7056;
    wire tmp7057;
    wire tmp7058;
    wire tmp7059;
    wire tmp7060;
    wire tmp7061;
    wire tmp7063;
    wire tmp7064;
    wire tmp7065;
    wire tmp7066;
    wire[7:0] tmp7079;
    wire tmp7080;
    wire[8:0] tmp7082;
    wire[8:0] tmp7093;
    wire[8:0] tmp7094;
    wire[9:0] tmp7097;
    wire tmp7098;
    wire tmp7099;
    wire tmp7100;
    wire tmp7101;
    wire tmp7103;
    wire tmp7104;
    wire tmp7105;
    wire tmp7106;
    wire tmp7107;
    wire tmp7109;
    wire[8:0] tmp7118;
    wire[8:0] tmp7119;
    wire[7:0] tmp7120;
    wire tmp7121;
    wire[8:0] tmp7123;
    wire tmp7125;
    wire tmp7126;
    wire[9:0] tmp7138;
    wire tmp7139;
    wire tmp7140;
    wire tmp7141;
    wire tmp7142;
    wire tmp7143;
    wire tmp7145;
    wire tmp7146;
    wire tmp7147;
    wire tmp7148;
    wire tmp7151;
    wire[8:0] tmp7157;
    wire[8:0] tmp7160;
    wire[7:0] tmp7161;
    wire tmp7162;
    wire[8:0] tmp7164;
    wire[8:0] tmp7176;
    wire[9:0] tmp7179;
    wire tmp7180;
    wire tmp7181;
    wire tmp7182;
    wire tmp7183;
    wire tmp7185;
    wire tmp7186;
    wire tmp7187;
    wire tmp7188;
    wire tmp7189;
    wire[6:0] tmp7226;
    wire tmp7227;
    wire[7:0] tmp7229;
    wire[6:0] tmp7249;
    wire tmp7250;
    wire[7:0] tmp7252;
    wire tmp7270;
    wire[6:0] tmp7272;
    wire tmp7273;
    wire[7:0] tmp7275;
    wire tmp7291;
    wire tmp7294;
    wire[6:0] tmp7295;
    wire tmp7296;
    wire[7:0] tmp7298;
    wire[7:0] tmp7319;
    wire[8:0] tmp7324;
    wire tmp7325;
    wire[8:0] tmp7336;
    wire tmp7340;
    wire tmp7343;
    wire tmp7344;
    wire tmp7350;
    wire tmp7353;
    wire tmp7356;
    wire tmp7365;
    wire tmp7368;
    wire tmp7369;
    wire tmp7370;
    wire tmp7371;
    wire tmp7385;
    wire tmp7390;
    wire tmp7393;
    wire[6:0] tmp7394;
    wire tmp7401;
    wire tmp7413;
    wire tmp7416;
    wire tmp7420;
    wire[8:0] tmp7425;
    wire tmp7426;
    wire[8:0] tmp7437;
    wire tmp7444;
    wire tmp7446;
    wire[7:0] tmp7449;
    wire[6:0] tmp7470;
    wire tmp7483;
    wire[8:0] tmp7488;
    wire tmp7489;
    wire tmp7492;
    wire tmp7495;
    wire tmp7496;
    wire tmp7508;
    wire tmp7520;
    wire tmp7523;
    wire[7:0] tmp7525;
    wire[6:0] tmp7546;
    wire[7:0] tmp7547;
    wire tmp7553;
    wire tmp7556;
    wire tmp7558;
    wire[8:0] tmp7564;
    wire tmp7565;
    wire tmp7567;
    wire tmp7568;
    wire tmp7571;
    wire tmp7572;
    wire tmp7579;
    wire tmp7581;
    wire tmp7584;
    wire[8:0] tmp7589;
    wire tmp7590;
    wire tmp7593;
    wire tmp7594;
    wire tmp7596;
    wire tmp7597;
    wire tmp7598;
    wire tmp7599;
    wire[7:0] tmp7600;
    wire[7:0] tmp7601;
    wire tmp7639;
    wire tmp7640;
    wire[7:0] tmp7692;
    wire[7:0] tmp7693;
    wire[7:0] tmp7694;
    wire[7:0] tmp7695;
    wire[7:0] tmp7696;
    wire[7:0] tmp7697;
    wire[7:0] tmp7698;
    wire[7:0] tmp7699;
    wire[7:0] tmp7700;
    wire[7:0] tmp7701;
    wire[7:0] tmp7702;
    wire[7:0] tmp7703;
    wire[7:0] tmp7704;
    wire[7:0] tmp7705;
    wire[7:0] tmp7706;
    wire[7:0] tmp7707;
    wire[7:0] tmp7708;
    wire[7:0] tmp7709;
    wire[7:0] tmp7710;
    wire[7:0] tmp7711;
    wire[7:0] tmp7712;
    wire[7:0] tmp7713;
    wire[7:0] tmp7714;
    wire[7:0] tmp7715;
    wire[7:0] tmp7716;
    wire[7:0] tmp7717;
    wire[7:0] tmp7718;
    wire[7:0] tmp7719;
    wire[7:0] tmp7720;
    wire[7:0] tmp7721;
    wire[7:0] tmp7722;
    wire[7:0] tmp7723;
    wire[7:0] tmp7724;
    wire[7:0] tmp7725;
    wire[7:0] tmp7726;
    wire[7:0] tmp7727;
    wire[7:0] tmp7728;
    wire[7:0] tmp7729;
    wire[7:0] tmp7730;
    wire[7:0] tmp7731;
    wire[7:0] tmp7732;
    wire[7:0] tmp7733;
    wire[7:0] tmp7734;
    wire[7:0] tmp7735;
    wire[7:0] tmp7736;
    wire[7:0] tmp7737;
    wire[7:0] tmp7738;
    wire[7:0] tmp7739;
    wire[7:0] tmp7740;
    wire[7:0] tmp7741;
    wire[7:0] tmp7742;
    wire[7:0] tmp7743;
    wire[7:0] tmp7744;
    wire[7:0] tmp7745;
    wire[7:0] tmp7746;
    wire[7:0] tmp7747;
    wire[7:0] tmp7748;
    wire[7:0] tmp7749;
    wire[7:0] tmp7750;
    wire[7:0] tmp7751;
    wire[7:0] tmp7752;
    wire[7:0] tmp7753;
    wire[7:0] tmp7754;
    wire[7:0] tmp7755;
    wire[7:0] tmp7756;
    wire[7:0] tmp7757;
    wire[7:0] tmp7758;
    wire[7:0] tmp7759;
    wire[7:0] tmp7760;
    wire[7:0] tmp7761;
    wire[7:0] tmp7762;
    wire[7:0] tmp7763;
    wire[7:0] tmp7764;
    wire[7:0] tmp7765;
    wire[7:0] tmp7766;
    wire[7:0] tmp7767;
    wire[7:0] tmp7768;
    wire[7:0] tmp7769;
    wire[7:0] tmp7770;
    wire[7:0] tmp7771;
    wire[7:0] tmp7772;
    wire[7:0] tmp7773;
    wire[7:0] tmp7774;
    wire[7:0] tmp7775;
    wire[7:0] tmp7776;
    wire[7:0] tmp7777;
    wire[7:0] tmp7778;
    wire[7:0] tmp7779;
    wire[7:0] tmp7780;
    wire[7:0] tmp7781;
    wire[7:0] tmp7782;
    wire[7:0] tmp7783;
    wire[7:0] tmp7784;
    wire[7:0] tmp7785;
    wire[7:0] tmp7786;
    wire[7:0] tmp7787;
    wire[7:0] tmp7788;
    wire[7:0] tmp7789;
    wire[7:0] tmp7790;
    wire[7:0] tmp7791;
    wire[7:0] tmp7792;
    wire[7:0] tmp7793;
    wire[7:0] tmp7794;
    wire[7:0] tmp7795;
    wire[7:0] tmp7796;
    wire[7:0] tmp7797;
    wire[7:0] tmp7798;
    wire[7:0] tmp7799;
    wire[7:0] tmp7800;
    wire[7:0] tmp7801;
    wire[7:0] tmp7802;
    wire[7:0] tmp7803;
    wire[7:0] tmp7804;
    wire[7:0] tmp7805;
    wire[7:0] tmp7806;
    wire[7:0] tmp7807;
    wire[7:0] tmp7808;
    wire[7:0] tmp7809;
    wire[7:0] tmp7810;
    wire[7:0] tmp7811;
    wire[7:0] tmp7812;
    wire[7:0] tmp7813;
    wire[7:0] tmp7814;
    wire[7:0] tmp7815;
    wire[7:0] tmp7816;
    wire[7:0] tmp7817;
    wire[7:0] tmp7818;
    wire[7:0] tmp7819;
    wire[7:0] tmp7820;
    wire[7:0] tmp7821;
    wire[7:0] tmp7822;
    wire[7:0] tmp7823;
    wire[7:0] tmp7824;
    wire[7:0] tmp7825;
    wire[7:0] tmp7826;
    wire[7:0] tmp7827;
    wire[7:0] tmp7828;
    wire[7:0] tmp7829;
    wire[7:0] tmp7830;
    wire[7:0] tmp7831;
    wire tmp7832;
    wire tmp7833;
    wire tmp7834;
    wire tmp7835;
    wire tmp7836;
    wire tmp7837;
    wire tmp7838;
    wire tmp7839;
    wire tmp7840;
    wire tmp7841;
    wire tmp7842;
    wire tmp7843;
    wire tmp7844;
    wire tmp7845;
    wire tmp7846;
    wire tmp7847;
    wire[3:0] tmp7848;
    wire[3:0] tmp7849;
    wire[3:0] tmp7850;
    wire[3:0] tmp7851;
    wire[3:0] tmp7852;
    wire[3:0] tmp7853;
    wire[3:0] tmp7854;
    wire[3:0] tmp7855;
    wire[3:0] tmp7856;
    wire[3:0] tmp7857;
    wire[3:0] tmp7858;
    wire[3:0] tmp7859;
    wire[3:0] tmp7860;
    wire[3:0] tmp7861;
    wire tmp7862;
    wire tmp7863;
    wire tmp7864;
    wire tmp7865;
    wire tmp7866;
    wire[7:0] tmp7869;
    wire[7:0] tmp7870;
    wire[7:0] tmp7873;
    wire[7:0] tmp7874;
    wire[7:0] tmp7877;
    wire[7:0] tmp7878;
    wire[7:0] tmp7881;
    wire[7:0] tmp7882;
    wire[7:0] tmp7885;
    wire[7:0] tmp7886;
    wire[7:0] tmp7889;
    wire[7:0] tmp7890;
    wire[7:0] tmp7893;
    wire[7:0] tmp7894;
    wire[7:0] tmp7897;
    wire[7:0] tmp7898;
    wire[2:0] tmp7903;
    wire[3:0] tmp7904;
    wire[3:0] tmp7905;
    wire tmp7908;
    wire tmp7914;
    wire tmp7917;
    wire tmp7918;
    wire tmp7919;
    wire tmp7920;
    wire tmp7921;
    wire tmp7923;
    wire[3:0] tmp7924;
    wire[4:0] tmp7925;
    wire[5:0] tmp7926;
    wire[4:0] tmp7927;
    wire[4:0] tmp7928;

    initial begin
        mem_0[0]=3'h4;
        mem_0[1]=3'h1;
        mem_0[2]=3'h2;
        mem_0[3]=3'h3;
        mem_0[4]=3'h1;
        mem_0[5]=3'h2;
        mem_0[6]=3'h3;
        mem_0[7]=3'h1;
        mem_0[8]=3'h2;
        mem_0[9]=3'h3;
        mem_0[10]=3'h1;
        mem_0[11]=3'h2;
        mem_0[12]=3'h3;
        mem_0[13]=3'h1;
        mem_0[14]=3'h2;
        mem_0[15]=3'h3;
        mem_0[16]=3'h1;
        mem_0[17]=3'h2;
        mem_0[18]=3'h3;
        mem_0[19]=3'h1;
        mem_0[20]=3'h2;
        mem_0[21]=3'h3;
        mem_0[22]=3'h1;
        mem_0[23]=3'h2;
        mem_0[24]=3'h3;
        mem_0[25]=3'h1;
        mem_0[26]=3'h2;
        mem_0[27]=3'h3;
        mem_0[28]=3'h1;
        mem_0[29]=3'h2;
        mem_0[30]=3'h3;
        mem_0[31]=3'h1;
    end

    initial begin
        mem_1[0]=4'h0;
        mem_1[1]=4'h4;
        mem_1[2]=4'h4;
        mem_1[3]=4'h4;
        mem_1[4]=4'hf;
        mem_1[5]=4'hf;
        mem_1[6]=4'hf;
        mem_1[7]=4'h0;
        mem_1[8]=4'h0;
        mem_1[9]=4'h0;
        mem_1[10]=4'h0;
        mem_1[11]=4'h0;
        mem_1[12]=4'h0;
        mem_1[13]=4'h0;
        mem_1[14]=4'h0;
        mem_1[15]=4'h0;
        mem_1[16]=4'h0;
        mem_1[17]=4'h0;
        mem_1[18]=4'h0;
        mem_1[19]=4'h0;
        mem_1[20]=4'h0;
        mem_1[21]=4'h0;
        mem_1[22]=4'h0;
        mem_1[23]=4'h0;
        mem_1[24]=4'h0;
        mem_1[25]=4'h0;
        mem_1[26]=4'h0;
        mem_1[27]=4'h0;
        mem_1[28]=4'h0;
        mem_1[29]=4'h0;
        mem_1[30]=4'h0;
        mem_1[31]=4'h0;
    end

    initial begin
        mem_2[0]=4'h0;
        mem_2[1]=4'h1;
        mem_2[2]=4'h1;
        mem_2[3]=4'h1;
        mem_2[4]=4'h4;
        mem_2[5]=4'h4;
        mem_2[6]=4'h4;
        mem_2[7]=4'hf;
        mem_2[8]=4'hf;
        mem_2[9]=4'hf;
        mem_2[10]=4'h0;
        mem_2[11]=4'h0;
        mem_2[12]=4'h0;
        mem_2[13]=4'h0;
        mem_2[14]=4'h0;
        mem_2[15]=4'h0;
        mem_2[16]=4'h0;
        mem_2[17]=4'h0;
        mem_2[18]=4'h0;
        mem_2[19]=4'h0;
        mem_2[20]=4'h0;
        mem_2[21]=4'h0;
        mem_2[22]=4'h0;
        mem_2[23]=4'h0;
        mem_2[24]=4'h0;
        mem_2[25]=4'h0;
        mem_2[26]=4'h0;
        mem_2[27]=4'h0;
        mem_2[28]=4'h0;
        mem_2[29]=4'h0;
        mem_2[30]=4'h0;
        mem_2[31]=4'h0;
    end

    // Combinational
    assign _ver_out_tmp_0 = 128;
    assign _ver_out_tmp_1 = 128;
    assign _ver_out_tmp_2 = 128;
    assign _ver_out_tmp_3 = 128;
    assign _ver_out_tmp_4 = 128;
    assign _ver_out_tmp_5 = 128;
    assign _ver_out_tmp_6 = 128;
    assign _ver_out_tmp_7 = 128;
    assign _ver_out_tmp_8 = 128;
    assign _ver_out_tmp_9 = 128;
    assign _ver_out_tmp_10 = 128;
    assign _ver_out_tmp_11 = 128;
    assign _ver_out_tmp_12 = 128;
    assign _ver_out_tmp_13 = 128;
    assign _ver_out_tmp_14 = 128;
    assign _ver_out_tmp_15 = 128;
    assign _ver_out_tmp_16 = 128;
    assign _ver_out_tmp_17 = 128;
    assign _ver_out_tmp_18 = 128;
    assign _ver_out_tmp_19 = 128;
    assign _ver_out_tmp_20 = 128;
    assign _ver_out_tmp_21 = 128;
    assign _ver_out_tmp_22 = 128;
    assign _ver_out_tmp_23 = 128;
    assign _ver_out_tmp_24 = 128;
    assign _ver_out_tmp_25 = 128;
    assign _ver_out_tmp_26 = 128;
    assign _ver_out_tmp_27 = 128;
    assign _ver_out_tmp_28 = 128;
    assign _ver_out_tmp_29 = 128;
    assign _ver_out_tmp_30 = 128;
    assign _ver_out_tmp_31 = 128;
    assign _ver_out_tmp_32 = 128;
    assign _ver_out_tmp_33 = 128;
    assign _ver_out_tmp_34 = 128;
    assign _ver_out_tmp_35 = 128;
    assign _ver_out_tmp_36 = 128;
    assign _ver_out_tmp_37 = 128;
    assign _ver_out_tmp_38 = 128;
    assign _ver_out_tmp_39 = 128;
    assign _ver_out_tmp_40 = 128;
    assign _ver_out_tmp_41 = 128;
    assign _ver_out_tmp_42 = 128;
    assign _ver_out_tmp_43 = 128;
    assign _ver_out_tmp_44 = 128;
    assign _ver_out_tmp_45 = 128;
    assign _ver_out_tmp_46 = 128;
    assign _ver_out_tmp_47 = 128;
    assign _ver_out_tmp_48 = 128;
    assign _ver_out_tmp_49 = 128;
    assign _ver_out_tmp_50 = 128;
    assign _ver_out_tmp_51 = 128;
    assign _ver_out_tmp_52 = 128;
    assign _ver_out_tmp_53 = 128;
    assign _ver_out_tmp_54 = 128;
    assign _ver_out_tmp_55 = 128;
    assign _ver_out_tmp_56 = 128;
    assign _ver_out_tmp_57 = 128;
    assign _ver_out_tmp_58 = 128;
    assign _ver_out_tmp_59 = 128;
    assign _ver_out_tmp_60 = 128;
    assign _ver_out_tmp_61 = 128;
    assign _ver_out_tmp_62 = 128;
    assign _ver_out_tmp_63 = 128;
    assign _ver_out_tmp_64 = 128;
    assign _ver_out_tmp_65 = 128;
    assign _ver_out_tmp_66 = 128;
    assign _ver_out_tmp_67 = 128;
    assign _ver_out_tmp_68 = 128;
    assign _ver_out_tmp_69 = 128;
    assign _ver_out_tmp_70 = 128;
    assign _ver_out_tmp_71 = 128;
    assign _ver_out_tmp_72 = 128;
    assign _ver_out_tmp_73 = 128;
    assign _ver_out_tmp_74 = 128;
    assign _ver_out_tmp_75 = 128;
    assign _ver_out_tmp_76 = 128;
    assign _ver_out_tmp_77 = 128;
    assign _ver_out_tmp_78 = 128;
    assign _ver_out_tmp_79 = 128;
    assign _ver_out_tmp_80 = 128;
    assign _ver_out_tmp_81 = 128;
    assign _ver_out_tmp_82 = 128;
    assign _ver_out_tmp_83 = 128;
    assign _ver_out_tmp_84 = 128;
    assign _ver_out_tmp_85 = 128;
    assign _ver_out_tmp_86 = 128;
    assign _ver_out_tmp_87 = 128;
    assign _ver_out_tmp_88 = 128;
    assign _ver_out_tmp_89 = 128;
    assign _ver_out_tmp_90 = 128;
    assign _ver_out_tmp_91 = 128;
    assign const_1_1 = 1;
    assign const_2_0 = 0;
    assign const_3_0 = 0;
    assign const_4_0 = 0;
    assign const_5_4 = 4;
    assign const_6_0 = 0;
    assign const_7_2 = 2;
    assign const_8_1 = 1;
    assign const_9_0 = 0;
    assign const_10_0 = 0;
    assign const_11_0 = 0;
    assign const_12_0 = 0;
    assign const_13_1 = 1;
    assign const_14_0 = 0;
    assign const_15_0 = 0;
    assign const_16_1 = 1;
    assign const_17_0 = 0;
    assign const_18_0 = 0;
    assign const_19_0 = 0;
    assign const_20_15 = 15;
    assign const_21_1 = 1;
    assign const_22_0 = 0;
    assign const_23_2 = 2;
    assign const_24_0 = 0;
    assign const_25_3 = 3;
    assign const_26_0 = 0;
    assign const_27_0 = 0;
    assign const_28_0 = 0;
    assign const_29_0 = 0;
    assign const_30_0 = 0;
    assign const_31_0 = 0;
    assign const_32_127 = 127;
    assign const_34_0 = 0;
    assign const_35_0 = 0;
    assign const_36_0 = 0;
    assign const_37_0 = 0;
    assign const_38_0 = 0;
    assign const_39_127 = 127;
    assign const_41_0 = 0;
    assign const_42_0 = 0;
    assign const_43_0 = 0;
    assign const_44_0 = 0;
    assign const_45_0 = 0;
    assign const_46_127 = 127;
    assign const_48_0 = 0;
    assign const_49_0 = 0;
    assign const_50_0 = 0;
    assign const_51_0 = 0;
    assign const_52_0 = 0;
    assign const_53_127 = 127;
    assign const_55_6 = 6;
    assign const_56_0 = 0;
    assign const_57_7 = 7;
    assign const_58_0 = 0;
    assign const_59_4 = 4;
    assign const_60_0 = 0;
    assign const_61_5 = 5;
    assign const_62_0 = 0;
    assign const_63_0 = 0;
    assign const_64_0 = 0;
    assign const_65_0 = 0;
    assign const_66_0 = 0;
    assign const_67_0 = 0;
    assign const_68_0 = 0;
    assign const_69_127 = 127;
    assign const_71_0 = 0;
    assign const_72_0 = 0;
    assign const_73_0 = 0;
    assign const_74_0 = 0;
    assign const_75_0 = 0;
    assign const_76_0 = 0;
    assign const_77_127 = 127;
    assign const_79_0 = 0;
    assign const_80_0 = 0;
    assign const_81_0 = 0;
    assign const_82_0 = 0;
    assign const_83_0 = 0;
    assign const_84_0 = 0;
    assign const_85_127 = 127;
    assign const_87_0 = 0;
    assign const_88_0 = 0;
    assign const_89_0 = 0;
    assign const_90_0 = 0;
    assign const_91_0 = 0;
    assign const_92_0 = 0;
    assign const_93_127 = 127;
    assign const_95_8 = 8;
    assign const_97_0 = 0;
    assign const_98_0 = 0;
    assign const_99_127 = 127;
    assign const_100_0 = 0;
    assign const_102_0 = 0;
    assign const_103_0 = 0;
    assign const_104_127 = 127;
    assign const_105_0 = 0;
    assign const_107_0 = 0;
    assign const_108_0 = 0;
    assign const_109_127 = 127;
    assign const_110_0 = 0;
    assign const_112_0 = 0;
    assign const_113_0 = 0;
    assign const_114_127 = 127;
    assign const_115_0 = 0;
    assign const_116_2 = 2;
    assign const_117_0 = 0;
    assign const_118_0 = 0;
    assign const_119_0 = 0;
    assign const_120_15 = 15;
    assign const_121_1 = 1;
    assign const_122_0 = 0;
    assign const_123_2 = 2;
    assign const_124_0 = 0;
    assign const_125_3 = 3;
    assign const_126_0 = 0;
    assign const_127_0 = 0;
    assign const_128_0 = 0;
    assign const_129_0 = 0;
    assign const_130_0 = 0;
    assign const_131_0 = 0;
    assign const_132_127 = 127;
    assign const_134_0 = 0;
    assign const_135_0 = 0;
    assign const_136_0 = 0;
    assign const_137_0 = 0;
    assign const_138_0 = 0;
    assign const_139_127 = 127;
    assign const_141_0 = 0;
    assign const_142_0 = 0;
    assign const_143_0 = 0;
    assign const_144_0 = 0;
    assign const_145_0 = 0;
    assign const_146_127 = 127;
    assign const_148_0 = 0;
    assign const_149_0 = 0;
    assign const_150_0 = 0;
    assign const_151_0 = 0;
    assign const_152_0 = 0;
    assign const_153_127 = 127;
    assign const_155_6 = 6;
    assign const_156_0 = 0;
    assign const_157_7 = 7;
    assign const_158_0 = 0;
    assign const_159_4 = 4;
    assign const_160_0 = 0;
    assign const_161_5 = 5;
    assign const_162_0 = 0;
    assign const_163_0 = 0;
    assign const_164_0 = 0;
    assign const_165_0 = 0;
    assign const_166_0 = 0;
    assign const_167_0 = 0;
    assign const_168_0 = 0;
    assign const_169_127 = 127;
    assign const_171_0 = 0;
    assign const_172_0 = 0;
    assign const_173_0 = 0;
    assign const_174_0 = 0;
    assign const_175_0 = 0;
    assign const_176_0 = 0;
    assign const_177_127 = 127;
    assign const_179_0 = 0;
    assign const_180_0 = 0;
    assign const_181_0 = 0;
    assign const_182_0 = 0;
    assign const_183_0 = 0;
    assign const_184_0 = 0;
    assign const_185_127 = 127;
    assign const_187_0 = 0;
    assign const_188_0 = 0;
    assign const_189_0 = 0;
    assign const_190_0 = 0;
    assign const_191_0 = 0;
    assign const_192_0 = 0;
    assign const_193_127 = 127;
    assign const_195_8 = 8;
    assign const_197_0 = 0;
    assign const_198_0 = 0;
    assign const_199_127 = 127;
    assign const_200_0 = 0;
    assign const_202_0 = 0;
    assign const_203_0 = 0;
    assign const_204_127 = 127;
    assign const_205_0 = 0;
    assign const_207_0 = 0;
    assign const_208_0 = 0;
    assign const_209_127 = 127;
    assign const_210_0 = 0;
    assign const_212_0 = 0;
    assign const_213_0 = 0;
    assign const_214_127 = 127;
    assign const_215_0 = 0;
    assign const_216_3 = 3;
    assign const_217_0 = 0;
    assign const_218_0 = 0;
    assign const_219_0 = 0;
    assign const_220_0 = 0;
    assign const_221_0 = 0;
    assign const_222_0 = 0;
    assign const_223_0 = 0;
    assign const_224_0 = 0;
    assign const_225_0 = 0;
    assign const_226_0 = 0;
    assign const_227_0 = 0;
    assign const_228_0 = 0;
    assign const_229_0 = 0;
    assign const_230_0 = 0;
    assign const_231_0 = 0;
    assign const_232_0 = 0;
    assign const_233_0 = 0;
    assign const_234_0 = 0;
    assign const_235_0 = 0;
    assign const_236_0 = 0;
    assign const_237_0 = 0;
    assign const_238_0 = 0;
    assign const_239_0 = 0;
    assign const_241_0 = 0;
    assign const_242_0 = 0;
    assign const_243_127 = 127;
    assign const_244_0 = 0;
    assign const_246_0 = 0;
    assign const_247_0 = 0;
    assign const_248_127 = 127;
    assign const_249_0 = 0;
    assign const_251_0 = 0;
    assign const_252_0 = 0;
    assign const_253_127 = 127;
    assign const_254_0 = 0;
    assign const_256_0 = 0;
    assign const_257_0 = 0;
    assign const_258_127 = 127;
    assign const_259_0 = 0;
    assign const_261_0 = 0;
    assign const_262_0 = 0;
    assign const_263_127 = 127;
    assign const_264_0 = 0;
    assign const_266_0 = 0;
    assign const_267_0 = 0;
    assign const_268_127 = 127;
    assign const_269_0 = 0;
    assign const_271_0 = 0;
    assign const_272_0 = 0;
    assign const_273_127 = 127;
    assign const_274_0 = 0;
    assign const_276_0 = 0;
    assign const_277_0 = 0;
    assign const_278_127 = 127;
    assign const_279_0 = 0;
    assign const_280_0 = 0;
    assign const_281_0 = 0;
    assign const_282_0 = 0;
    assign const_283_0 = 0;
    assign const_284_0 = 0;
    assign const_285_0 = 0;
    assign const_286_0 = 0;
    assign const_287_0 = 0;
    assign const_288_0 = 0;
    assign const_289_0 = 0;
    assign const_290_15 = 15;
    assign const_291_0 = 0;
    assign const_292_0 = 0;
    assign const_293_0 = 0;
    assign const_294_8 = 8;
    assign const_295_0 = 0;
    assign const_297_0 = 0;
    assign const_298_0 = 0;
    assign const_299_127 = 127;
    assign const_300_0 = 0;
    assign const_302_0 = 0;
    assign const_303_0 = 0;
    assign const_304_127 = 127;
    assign const_305_0 = 0;
    assign const_307_0 = 0;
    assign const_308_0 = 0;
    assign const_309_127 = 127;
    assign const_310_0 = 0;
    assign const_312_0 = 0;
    assign const_313_0 = 0;
    assign const_314_127 = 127;
    assign const_315_0 = 0;
    assign const_316_1 = 1;
    assign const_317_0 = 0;
    assign const_318_0 = 0;
    assign const_319_0 = 0;
    assign const_320_0 = 0;
    assign const_321_0 = 0;
    assign const_322_0 = 0;
    assign const_323_127 = 127;
    assign const_325_0 = 0;
    assign const_326_0 = 0;
    assign const_327_0 = 0;
    assign const_328_0 = 0;
    assign const_329_0 = 0;
    assign const_330_127 = 127;
    assign const_332_0 = 0;
    assign const_333_0 = 0;
    assign const_334_0 = 0;
    assign const_335_0 = 0;
    assign const_336_0 = 0;
    assign const_337_127 = 127;
    assign const_339_0 = 0;
    assign const_340_0 = 0;
    assign const_341_0 = 0;
    assign const_342_0 = 0;
    assign const_343_0 = 0;
    assign const_344_127 = 127;
    assign const_346_4 = 4;
    assign const_347_0 = 0;
    assign const_349_0 = 0;
    assign const_350_0 = 0;
    assign const_351_127 = 127;
    assign const_352_0 = 0;
    assign const_353_0 = 0;
    assign const_354_0 = 0;
    assign const_355_0 = 0;
    assign const_356_0 = 0;
    assign const_357_0 = 0;
    assign const_358_0 = 0;
    assign const_359_127 = 127;
    assign const_362_0 = 0;
    assign const_363_0 = 0;
    assign const_364_127 = 127;
    assign const_365_0 = 0;
    assign const_366_0 = 0;
    assign const_367_0 = 0;
    assign const_368_0 = 0;
    assign const_369_0 = 0;
    assign const_370_0 = 0;
    assign const_371_0 = 0;
    assign const_372_127 = 127;
    assign const_375_0 = 0;
    assign const_376_0 = 0;
    assign const_377_127 = 127;
    assign const_378_0 = 0;
    assign const_379_0 = 0;
    assign const_380_0 = 0;
    assign const_381_0 = 0;
    assign const_382_0 = 0;
    assign const_383_0 = 0;
    assign const_384_0 = 0;
    assign const_385_127 = 127;
    assign const_388_0 = 0;
    assign const_389_0 = 0;
    assign const_390_127 = 127;
    assign const_391_0 = 0;
    assign const_392_0 = 0;
    assign const_393_0 = 0;
    assign const_394_0 = 0;
    assign const_395_0 = 0;
    assign const_396_0 = 0;
    assign const_397_0 = 0;
    assign const_398_127 = 127;
    assign const_400_6 = 6;
    assign const_401_0 = 0;
    assign const_402_0 = 0;
    assign const_403_0 = 0;
    assign const_404_0 = 0;
    assign const_405_0 = 0;
    assign const_406_0 = 0;
    assign const_407_127 = 127;
    assign const_409_0 = 0;
    assign const_410_0 = 0;
    assign const_411_0 = 0;
    assign const_412_0 = 0;
    assign const_413_0 = 0;
    assign const_414_127 = 127;
    assign const_416_0 = 0;
    assign const_417_0 = 0;
    assign const_418_0 = 0;
    assign const_419_0 = 0;
    assign const_420_0 = 0;
    assign const_421_127 = 127;
    assign const_423_0 = 0;
    assign const_424_0 = 0;
    assign const_425_0 = 0;
    assign const_426_0 = 0;
    assign const_427_0 = 0;
    assign const_428_127 = 127;
    assign const_430_2 = 2;
    assign const_431_0 = 0;
    assign const_432_0 = 0;
    assign const_433_0 = 0;
    assign const_434_0 = 0;
    assign const_435_0 = 0;
    assign const_436_0 = 0;
    assign const_437_127 = 127;
    assign const_439_0 = 0;
    assign const_440_0 = 0;
    assign const_441_0 = 0;
    assign const_442_0 = 0;
    assign const_443_0 = 0;
    assign const_444_127 = 127;
    assign const_446_0 = 0;
    assign const_447_0 = 0;
    assign const_448_0 = 0;
    assign const_449_0 = 0;
    assign const_450_0 = 0;
    assign const_451_127 = 127;
    assign const_453_0 = 0;
    assign const_454_0 = 0;
    assign const_455_0 = 0;
    assign const_456_0 = 0;
    assign const_457_0 = 0;
    assign const_458_127 = 127;
    assign const_460_0 = 0;
    assign const_461_0 = 0;
    assign const_462_0 = 0;
    assign const_463_0 = 0;
    assign const_464_0 = 0;
    assign const_465_127 = 127;
    assign const_467_0 = 0;
    assign const_468_0 = 0;
    assign const_469_0 = 0;
    assign const_470_0 = 0;
    assign const_471_0 = 0;
    assign const_472_127 = 127;
    assign const_474_0 = 0;
    assign const_475_0 = 0;
    assign const_476_0 = 0;
    assign const_477_0 = 0;
    assign const_478_0 = 0;
    assign const_479_127 = 127;
    assign const_481_0 = 0;
    assign const_482_0 = 0;
    assign const_483_0 = 0;
    assign const_484_0 = 0;
    assign const_485_0 = 0;
    assign const_486_127 = 127;
    assign const_488_0 = 0;
    assign const_489_0 = 0;
    assign const_490_0 = 0;
    assign const_491_0 = 0;
    assign const_492_0 = 0;
    assign const_493_127 = 127;
    assign const_495_0 = 0;
    assign const_496_0 = 0;
    assign const_497_0 = 0;
    assign const_498_0 = 0;
    assign const_499_0 = 0;
    assign const_500_127 = 127;
    assign const_502_0 = 0;
    assign const_503_0 = 0;
    assign const_504_0 = 0;
    assign const_505_0 = 0;
    assign const_506_0 = 0;
    assign const_507_127 = 127;
    assign const_509_0 = 0;
    assign const_510_0 = 0;
    assign const_511_0 = 0;
    assign const_512_0 = 0;
    assign const_513_0 = 0;
    assign const_514_127 = 127;
    assign const_516_5 = 5;
    assign const_517_1 = 1;
    assign const_519_0 = 0;
    assign const_520_0 = 0;
    assign const_521_127 = 127;
    assign const_522_0 = 0;
    assign const_523_0 = 0;
    assign const_524_0 = 0;
    assign const_525_0 = 0;
    assign const_526_0 = 0;
    assign const_527_0 = 0;
    assign const_528_0 = 0;
    assign const_529_127 = 127;
    assign const_532_0 = 0;
    assign const_533_0 = 0;
    assign const_534_127 = 127;
    assign const_535_0 = 0;
    assign const_536_0 = 0;
    assign const_537_0 = 0;
    assign const_538_0 = 0;
    assign const_539_0 = 0;
    assign const_540_0 = 0;
    assign const_541_0 = 0;
    assign const_542_127 = 127;
    assign const_545_0 = 0;
    assign const_546_0 = 0;
    assign const_547_127 = 127;
    assign const_548_0 = 0;
    assign const_549_0 = 0;
    assign const_550_0 = 0;
    assign const_551_0 = 0;
    assign const_552_0 = 0;
    assign const_553_0 = 0;
    assign const_554_0 = 0;
    assign const_555_127 = 127;
    assign const_558_0 = 0;
    assign const_559_0 = 0;
    assign const_560_127 = 127;
    assign const_561_0 = 0;
    assign const_562_0 = 0;
    assign const_563_0 = 0;
    assign const_564_0 = 0;
    assign const_565_0 = 0;
    assign const_566_0 = 0;
    assign const_567_0 = 0;
    assign const_568_127 = 127;
    assign const_570_0 = 0;
    assign const_571_0 = 0;
    assign const_572_0 = 0;
    assign const_573_0 = 0;
    assign const_574_1 = 1;
    assign const_576_0 = 0;
    assign const_577_0 = 0;
    assign const_578_127 = 127;
    assign const_579_0 = 0;
    assign const_580_0 = 0;
    assign const_581_1 = 1;
    assign const_583_0 = 0;
    assign const_584_0 = 0;
    assign const_585_127 = 127;
    assign const_586_0 = 0;
    assign const_587_0 = 0;
    assign const_588_1 = 1;
    assign const_590_0 = 0;
    assign const_591_0 = 0;
    assign const_592_127 = 127;
    assign const_593_0 = 0;
    assign const_594_0 = 0;
    assign const_595_1 = 1;
    assign const_597_0 = 0;
    assign const_598_0 = 0;
    assign const_599_127 = 127;
    assign const_600_0 = 0;
    assign const_601_0 = 0;
    assign const_602_1 = 1;
    assign const_604_0 = 0;
    assign const_605_0 = 0;
    assign const_606_127 = 127;
    assign const_607_0 = 0;
    assign const_608_0 = 0;
    assign const_609_1 = 1;
    assign const_611_0 = 0;
    assign const_612_0 = 0;
    assign const_613_127 = 127;
    assign const_614_0 = 0;
    assign const_615_0 = 0;
    assign const_616_1 = 1;
    assign const_618_0 = 0;
    assign const_619_0 = 0;
    assign const_620_127 = 127;
    assign const_621_0 = 0;
    assign const_622_0 = 0;
    assign const_623_1 = 1;
    assign const_625_0 = 0;
    assign const_626_0 = 0;
    assign const_627_127 = 127;
    assign const_628_0 = 0;
    assign const_629_0 = 0;
    assign const_630_7 = 7;
    assign const_631_1 = 1;
    assign const_632_1 = 1;
    assign const_634_0 = 0;
    assign const_635_0 = 0;
    assign const_636_127 = 127;
    assign const_637_0 = 0;
    assign const_638_0 = 0;
    assign const_639_1 = 1;
    assign const_641_0 = 0;
    assign const_642_0 = 0;
    assign const_643_127 = 127;
    assign const_644_0 = 0;
    assign const_645_0 = 0;
    assign const_646_1 = 1;
    assign const_648_0 = 0;
    assign const_649_0 = 0;
    assign const_650_127 = 127;
    assign const_651_0 = 0;
    assign const_652_0 = 0;
    assign const_653_1 = 1;
    assign const_655_0 = 0;
    assign const_656_0 = 0;
    assign const_657_127 = 127;
    assign const_658_0 = 0;
    assign const_659_0 = 0;
    assign const_660_1 = 1;
    assign const_662_0 = 0;
    assign const_663_0 = 0;
    assign const_664_127 = 127;
    assign const_665_0 = 0;
    assign const_666_0 = 0;
    assign const_667_1 = 1;
    assign const_669_0 = 0;
    assign const_670_0 = 0;
    assign const_671_127 = 127;
    assign const_672_0 = 0;
    assign const_673_0 = 0;
    assign const_674_1 = 1;
    assign const_676_0 = 0;
    assign const_677_0 = 0;
    assign const_678_127 = 127;
    assign const_679_0 = 0;
    assign const_680_0 = 0;
    assign const_681_1 = 1;
    assign const_683_0 = 0;
    assign const_684_0 = 0;
    assign const_685_127 = 127;
    assign const_686_0 = 0;
    assign const_687_0 = 0;
    assign const_688_3 = 3;
    assign const_689_1 = 1;
    assign const_690_0 = 0;
    assign const_691_0 = 0;
    assign const_692_0 = 0;
    assign const_693_0 = 0;
    assign const_694_0 = 0;
    assign const_695_127 = 127;
    assign const_697_0 = 0;
    assign const_698_0 = 0;
    assign const_699_0 = 0;
    assign const_700_0 = 0;
    assign const_701_0 = 0;
    assign const_702_127 = 127;
    assign const_704_0 = 0;
    assign const_705_0 = 0;
    assign const_706_0 = 0;
    assign const_707_0 = 0;
    assign const_708_0 = 0;
    assign const_709_127 = 127;
    assign const_711_0 = 0;
    assign const_712_0 = 0;
    assign const_713_0 = 0;
    assign const_714_0 = 0;
    assign const_715_0 = 0;
    assign const_716_127 = 127;
    assign const_718_0 = 0;
    assign const_719_0 = 0;
    assign const_720_0 = 0;
    assign const_721_0 = 0;
    assign const_722_0 = 0;
    assign const_723_0 = 0;
    assign const_724_0 = 0;
    assign const_725_0 = 0;
    assign const_726_0 = 0;
    assign const_727_0 = 0;
    assign const_728_0 = 0;
    assign const_729_0 = 0;
    assign const_730_0 = 0;
    assign const_731_0 = 0;
    assign const_732_0 = 0;
    assign const_733_0 = 0;
    assign const_734_0 = 0;
    assign const_735_0 = 0;
    assign const_736_0 = 0;
    assign const_737_0 = 0;
    assign const_738_0 = 0;
    assign const_739_0 = 0;
    assign const_740_0 = 0;
    assign const_741_0 = 0;
    assign const_742_0 = 0;
    assign const_743_1 = 1;
    assign const_744_0 = 0;
    assign const_745_1 = 1;
    assign const_746_0 = 0;
    assign const_747_4 = 4;
    assign const_748_0 = 0;
    assign const_749_15 = 15;
    assign const_750_1 = 1;
    assign const_751_0 = 0;
    assign const_756_0 = 0;
    assign const_757_0 = 0;
    assign const_758_0 = 0;
    assign const_759_0 = 0;
    assign blue_o = tmp7920;
    assign green_o = tmp7914;
    assign red_o = tmp7908;
    assign tmp1 = {const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0};
    assign tmp2 = {tmp1, const_1_1};
    assign tmp3 = tmp0 + tmp2;
    assign tmp4 = {tmp3[26], tmp3[25], tmp3[24], tmp3[23], tmp3[22], tmp3[21], tmp3[20], tmp3[19], tmp3[18], tmp3[17], tmp3[16], tmp3[15], tmp3[14], tmp3[13], tmp3[12], tmp3[11], tmp3[10], tmp3[9], tmp3[8], tmp3[7], tmp3[6], tmp3[5], tmp3[4], tmp3[3], tmp3[2], tmp3[1], tmp3[0]};
    assign tmp8 = tmp5 == tmp7921;
    assign tmp32 = ~was_toggled;
    assign tmp34 = {tmp133, const_3_0};
    assign tmp35 = my_calculator_ctrl == tmp34;
    assign tmp36 = my_calculator_ctrl == const_5_4;
    assign tmp68 = tmp858 & tmp36;
    assign tmp78 = {tmp133, const_16_1};
    assign tmp79 = my_calculator_ctrl == tmp78;
    assign tmp87 = {tmp126, const_18_0};
    assign tmp88 = my_calculator_in_x == tmp87;
    assign tmp89 = my_calculator_in_x == const_20_15;
    assign tmp107 = tmp999 & tmp89;
    assign tmp126 = {const_22_0, const_22_0, const_22_0};
    assign tmp127 = {tmp126, const_21_1};
    assign tmp128 = my_calculator_in_x == tmp127;
    assign tmp130 = {tmp133, const_23_2};
    assign tmp131 = my_calculator_in_x == tmp130;
    assign tmp132 = tmp128 | tmp131;
    assign tmp133 = {const_26_0, const_26_0};
    assign tmp135 = my_calculator_in_x == tmp1175;
    assign tmp136 = tmp132 | tmp135;
    assign tmp137 = {tmp10[6], tmp10[5], tmp10[4], tmp10[3], tmp10[2], tmp10[1], tmp10[0]};
    assign tmp138 = {tmp137, const_27_0};
    assign tmp155 = tmp138 - tmp5375;
    assign tmp156 = {tmp155[8]};
    assign tmp157 = {tmp138[7]};
    assign tmp159 = tmp156 ^ tmp1227;
    assign tmp162 = tmp159 ^ tmp1604;
    assign tmp190 = tmp2787 & tmp1230;
    assign tmp192 = tmp190 ? _ver_out_tmp_44 : tmp1232;
    assign tmp204 = {tmp11[6], tmp11[5], tmp11[4], tmp11[3], tmp11[2], tmp11[1], tmp11[0]};
    assign tmp205 = {tmp204, const_34_0};
    assign tmp211 = {tmp657[8]};
    assign tmp216 = ~tmp6761;
    assign tmp217 = tmp661 ^ tmp216;
    assign tmp222 = tmp205 - tmp5375;
    assign tmp223 = {tmp222[8]};
    assign tmp224 = {tmp205[7]};
    assign tmp226 = tmp223 ^ tmp253;
    assign tmp229 = tmp226 ^ tmp1604;
    assign tmp230 = tmp217 & tmp229;
    assign tmp247 = tmp5375 - tmp205;
    assign tmp248 = {tmp247[8]};
    assign tmp251 = tmp248 ^ tmp1604;
    assign tmp253 = ~tmp224;
    assign tmp254 = tmp251 ^ tmp253;
    assign tmp255 = tmp5375 == tmp205;
    assign tmp256 = tmp254 | tmp255;
    assign tmp257 = tmp2236 & tmp256;
    assign tmp258 = tmp230 ? const_39_127 : tmp205;
    assign tmp259 = tmp257 ? _ver_out_tmp_84 : tmp258;
    assign tmp266 = ~tmp88;
    assign tmp281 = tmp7325 ^ tmp1604;
    assign tmp283 = ~tmp1893;
    assign tmp314 = tmp5375 - tmp7319;
    assign tmp320 = ~tmp1336;
    assign tmp325 = tmp7344 ? const_46_127 : tmp7319;
    assign tmp326 = tmp7371 ? _ver_out_tmp_49 : tmp325;
    assign tmp337 = tmp1025 & tmp136;
    assign tmp339 = {tmp7394, const_48_0};
    assign tmp344 = tmp5375 - tmp15;
    assign tmp348 = tmp7401 ^ tmp1604;
    assign tmp349 = {tmp15[7]};
    assign tmp356 = tmp339 - tmp5375;
    assign tmp358 = {tmp339[7]};
    assign tmp359 = ~tmp358;
    assign tmp363 = tmp7416 ^ tmp1604;
    assign tmp382 = {tmp7437[8]};
    assign tmp385 = tmp382 ^ tmp1604;
    assign tmp389 = tmp5375 == tmp339;
    assign tmp391 = tmp2323 & tmp7446;
    assign tmp392 = tmp7420 ? const_53_127 : tmp339;
    assign tmp407 = my_calculator_in_x == tmp1455;
    assign tmp409 = {const_58_0, const_57_7};
    assign tmp410 = my_calculator_in_x == tmp409;
    assign tmp411 = tmp407 | tmp410;
    assign tmp422 = ~tmp136;
    assign tmp489 = tmp501 & tmp411;
    assign tmp501 = tmp1025 & tmp422;
    assign tmp517 = {const_60_0, const_59_4};
    assign tmp518 = my_calculator_in_x == tmp517;
    assign tmp521 = my_calculator_in_x == tmp1585;
    assign tmp522 = tmp518 | tmp521;
    assign tmp525 = {tmp7026, tmp10};
    assign tmp529 = tmp525 + tmp1715;
    assign tmp530 = {tmp529[8], tmp529[7], tmp529[6], tmp529[5], tmp529[4], tmp529[3], tmp529[2], tmp529[1], tmp529[0]};
    assign tmp531 = {tmp530[7], tmp530[6], tmp530[5], tmp530[4], tmp530[3], tmp530[2], tmp530[1], tmp530[0]};
    assign tmp537 = {tmp6732[8]};
    assign tmp542 = ~tmp7026;
    assign tmp543 = tmp1188 ^ tmp542;
    assign tmp548 = tmp5375 - tmp12;
    assign tmp549 = {tmp548[8]};
    assign tmp552 = tmp549 ^ tmp1604;
    assign tmp556 = tmp543 & tmp1260;
    assign tmp561 = tmp531 - tmp5375;
    assign tmp562 = {tmp561[8]};
    assign tmp563 = {tmp531[7]};
    assign tmp564 = ~tmp563;
    assign tmp565 = tmp562 ^ tmp564;
    assign tmp568 = tmp565 ^ tmp1604;
    assign tmp569 = tmp531 == tmp5375;
    assign tmp570 = tmp568 | tmp569;
    assign tmp571 = tmp556 & tmp570;
    assign tmp589 = {tmp1766[8]};
    assign tmp595 = tmp1770 ^ tmp1604;
    assign tmp596 = tmp2787 & tmp595;
    assign tmp601 = tmp5375 - tmp531;
    assign tmp602 = {tmp601[8]};
    assign tmp605 = tmp602 ^ tmp1604;
    assign tmp608 = tmp605 ^ tmp564;
    assign tmp610 = tmp608 | tmp569;
    assign tmp611 = tmp596 & tmp610;
    assign tmp612 = tmp571 ? const_69_127 : tmp531;
    assign tmp613 = tmp611 ? _ver_out_tmp_24 : tmp612;
    assign tmp646 = {tmp6761, tmp11};
    assign tmp649 = {tmp711, tmp13};
    assign tmp650 = tmp646 + tmp649;
    assign tmp651 = {tmp650[8], tmp650[7], tmp650[6], tmp650[5], tmp650[4], tmp650[3], tmp650[2], tmp650[1], tmp650[0]};
    assign tmp652 = {tmp651[7], tmp651[6], tmp651[5], tmp651[4], tmp651[3], tmp651[2], tmp651[1], tmp651[0]};
    assign tmp657 = tmp5375 - tmp11;
    assign tmp661 = tmp211 ^ tmp1604;
    assign tmp670 = {tmp2516[8]};
    assign tmp673 = tmp670 ^ tmp1604;
    assign tmp676 = tmp673 ^ tmp1781;
    assign tmp677 = tmp217 & tmp676;
    assign tmp682 = tmp652 - tmp5375;
    assign tmp683 = {tmp682[8]};
    assign tmp684 = {tmp652[7]};
    assign tmp686 = tmp683 ^ tmp728;
    assign tmp689 = tmp686 ^ tmp1604;
    assign tmp690 = tmp652 == tmp5375;
    assign tmp691 = tmp689 | tmp690;
    assign tmp692 = tmp677 & tmp691;
    assign tmp701 = tmp2230 ^ tmp216;
    assign tmp711 = {tmp13[7]};
    assign tmp713 = tmp1779 ^ tmp1781;
    assign tmp717 = tmp2236 & tmp2274;
    assign tmp722 = tmp5375 - tmp652;
    assign tmp723 = {tmp722[8]};
    assign tmp726 = tmp723 ^ tmp1604;
    assign tmp728 = ~tmp684;
    assign tmp729 = tmp726 ^ tmp728;
    assign tmp731 = tmp729 | tmp690;
    assign tmp732 = tmp717 & tmp731;
    assign tmp733 = tmp692 ? const_77_127 : tmp652;
    assign tmp734 = tmp732 ? _ver_out_tmp_64 : tmp733;
    assign tmp767 = {tmp1893, tmp14};
    assign tmp770 = {tmp1396, tmp16};
    assign tmp771 = tmp767 + tmp770;
    assign tmp772 = {tmp771[8], tmp771[7], tmp771[6], tmp771[5], tmp771[4], tmp771[3], tmp771[2], tmp771[1], tmp771[0]};
    assign tmp773 = {tmp772[7], tmp772[6], tmp772[5], tmp772[4], tmp772[3], tmp772[2], tmp772[1], tmp772[0]};
    assign tmp798 = tmp1858 & tmp7483;
    assign tmp803 = tmp773 - tmp5375;
    assign tmp804 = {tmp803[8]};
    assign tmp805 = {tmp773[7]};
    assign tmp806 = ~tmp805;
    assign tmp807 = tmp804 ^ tmp806;
    assign tmp810 = tmp807 ^ tmp1604;
    assign tmp811 = tmp773 == tmp5375;
    assign tmp812 = tmp810 | tmp811;
    assign tmp813 = tmp798 & tmp812;
    assign tmp830 = tmp16 - tmp5375;
    assign tmp831 = {tmp830[8]};
    assign tmp838 = tmp7356 & tmp7508;
    assign tmp843 = tmp5375 - tmp773;
    assign tmp844 = {tmp843[8]};
    assign tmp847 = tmp844 ^ tmp1604;
    assign tmp850 = tmp847 ^ tmp806;
    assign tmp852 = tmp850 | tmp811;
    assign tmp853 = tmp838 & tmp852;
    assign tmp854 = tmp813 ? const_85_127 : tmp773;
    assign tmp855 = tmp853 ? _ver_out_tmp_69 : tmp854;
    assign tmp858 = tmp1145 & tmp4798;
    assign tmp888 = {tmp349, tmp15};
    assign tmp892 = tmp888 + tmp1968;
    assign tmp893 = {tmp892[8], tmp892[7], tmp892[6], tmp892[5], tmp892[4], tmp892[3], tmp892[2], tmp892[1], tmp892[0]};
    assign tmp894 = {tmp893[7], tmp893[6], tmp893[5], tmp893[4], tmp893[3], tmp893[2], tmp893[1], tmp893[0]};
    assign tmp918 = tmp7556 ^ tmp7558;
    assign tmp919 = tmp1870 & tmp918;
    assign tmp924 = tmp894 - tmp5375;
    assign tmp925 = {tmp924[8]};
    assign tmp926 = {tmp894[7]};
    assign tmp927 = ~tmp926;
    assign tmp928 = tmp925 ^ tmp927;
    assign tmp931 = tmp928 ^ tmp1604;
    assign tmp933 = tmp931 | tmp972;
    assign tmp934 = tmp919 & tmp933;
    assign tmp942 = ~tmp349;
    assign tmp951 = tmp17 - tmp5375;
    assign tmp959 = tmp2323 & tmp7584;
    assign tmp964 = tmp5375 - tmp894;
    assign tmp965 = {tmp964[8]};
    assign tmp968 = tmp965 ^ tmp1604;
    assign tmp971 = tmp968 ^ tmp927;
    assign tmp972 = tmp5375 == tmp894;
    assign tmp973 = tmp971 | tmp972;
    assign tmp974 = tmp959 & tmp973;
    assign tmp975 = tmp934 ? const_93_127 : tmp894;
    assign tmp976 = tmp974 ? _ver_out_tmp_71 : tmp975;
    assign tmp997 = tmp1070 & tmp79;
    assign tmp999 = tmp997 & tmp266;
    assign tmp1000 = ~tmp89;
    assign tmp1006 = tmp1104 & tmp522;
    assign tmp1007 = my_calculator_in_x == const_95_8;
    assign tmp1015 = {tmp7034[7], tmp7034[6], tmp7034[5], tmp7034[4], tmp7034[3], tmp7034[2], tmp7034[1], tmp7034[0]};
    assign tmp1025 = tmp999 & tmp1000;
    assign tmp1030 = ~tmp522;
    assign tmp1056 = tmp1104 & tmp1030;
    assign tmp1064 = tmp2532 ? tmp4109 : tmp7324;
    assign tmp1070 = tmp858 & tmp5081;
    assign tmp1083 = tmp15 == _ver_out_tmp_83;
    assign tmp1089 = tmp1083 ? tmp4109 : tmp344;
    assign tmp1103 = ~tmp411;
    assign tmp1104 = tmp501 & tmp1103;
    assign tmp1107 = tmp1056 & tmp1007;
    assign tmp1109 = {const_117_0, const_116_2};
    assign tmp1110 = my_calculator_ctrl == tmp1109;
    assign tmp1121 = my_calculator_in_y == tmp87;
    assign tmp1122 = my_calculator_in_y == const_120_15;
    assign tmp1133 = tmp1545 & tmp1122;
    assign tmp1145 = ~tmp32;
    assign tmp1169 = my_calculator_in_y == tmp127;
    assign tmp1172 = my_calculator_in_y == tmp130;
    assign tmp1173 = tmp1169 | tmp1172;
    assign tmp1175 = {tmp133, const_125_3};
    assign tmp1176 = my_calculator_in_y == tmp1175;
    assign tmp1177 = tmp1173 | tmp1176;
    assign tmp1188 = tmp537 ^ tmp1604;
    assign tmp1204 = tmp543 & tmp162;
    assign tmp1221 = tmp5375 - tmp138;
    assign tmp1222 = {tmp1221[8]};
    assign tmp1225 = tmp1222 ^ tmp1604;
    assign tmp1227 = ~tmp157;
    assign tmp1228 = tmp1225 ^ tmp1227;
    assign tmp1229 = tmp5375 == tmp138;
    assign tmp1230 = tmp1228 | tmp1229;
    assign tmp1232 = tmp1204 ? const_132_127 : tmp138;
    assign tmp1247 = {tmp12[6], tmp12[5], tmp12[4], tmp12[3], tmp12[2], tmp12[1], tmp12[0]};
    assign tmp1248 = {tmp1247, const_134_0};
    assign tmp1260 = tmp552 ^ tmp2258;
    assign tmp1265 = tmp1248 - tmp5375;
    assign tmp1266 = {tmp1265[8]};
    assign tmp1269 = tmp1266 ^ tmp1296;
    assign tmp1272 = tmp1269 ^ tmp1604;
    assign tmp1273 = tmp1260 & tmp1272;
    assign tmp1290 = tmp5375 - tmp1248;
    assign tmp1291 = {tmp1290[8]};
    assign tmp1294 = tmp1291 ^ tmp1604;
    assign tmp1295 = {tmp1248[7]};
    assign tmp1296 = ~tmp1295;
    assign tmp1297 = tmp1294 ^ tmp1296;
    assign tmp1298 = tmp5375 == tmp1248;
    assign tmp1299 = tmp1297 | tmp1298;
    assign tmp1300 = tmp595 & tmp1299;
    assign tmp1301 = tmp1273 ? const_139_127 : tmp1248;
    assign tmp1302 = tmp1300 ? _ver_out_tmp_3 : tmp1301;
    assign tmp1316 = {tmp14[6], tmp14[5], tmp14[4], tmp14[3], tmp14[2], tmp14[1], tmp14[0]};
    assign tmp1335 = {tmp7336[8]};
    assign tmp1336 = {tmp7319[7]};
    assign tmp1360 = {tmp314[8]};
    assign tmp1384 = tmp1832 & tmp1177;
    assign tmp1386 = {tmp7470, const_148_0};
    assign tmp1392 = {tmp2573[8]};
    assign tmp1395 = tmp1392 ^ tmp1604;
    assign tmp1396 = {tmp16[7]};
    assign tmp1420 = tmp831 ^ tmp2019;
    assign tmp1428 = tmp5375 - tmp1386;
    assign tmp1429 = {tmp1428[8]};
    assign tmp1432 = tmp1429 ^ tmp1604;
    assign tmp1433 = {tmp1386[7]};
    assign tmp1434 = ~tmp1433;
    assign tmp1436 = tmp5375 == tmp1386;
    assign tmp1437 = tmp7520 | tmp1436;
    assign tmp1439 = tmp7496 ? const_153_127 : tmp1386;
    assign tmp1455 = {const_156_0, const_155_6};
    assign tmp1456 = my_calculator_in_y == tmp1455;
    assign tmp1459 = my_calculator_in_y == tmp409;
    assign tmp1460 = tmp1456 | tmp1459;
    assign tmp1545 = tmp1953 & tmp2132;
    assign tmp1580 = tmp1692 & tmp1460;
    assign tmp1583 = my_calculator_in_y == tmp517;
    assign tmp1585 = {const_162_0, const_161_5};
    assign tmp1586 = my_calculator_in_y == tmp1585;
    assign tmp1587 = tmp1583 | tmp1586;
    assign tmp1594 = tmp525 + tmp646;
    assign tmp1595 = {tmp1594[8], tmp1594[7], tmp1594[6], tmp1594[5], tmp1594[4], tmp1594[3], tmp1594[2], tmp1594[1], tmp1594[0]};
    assign tmp1596 = {tmp1595[7], tmp1595[6], tmp1595[5], tmp1595[4], tmp1595[3], tmp1595[2], tmp1595[1], tmp1595[0]};
    assign tmp1604 = ~tmp1783;
    assign tmp1621 = tmp543 & tmp217;
    assign tmp1626 = tmp1596 - tmp5375;
    assign tmp1627 = {tmp1626[8]};
    assign tmp1630 = tmp1627 ^ tmp1672;
    assign tmp1633 = tmp1630 ^ tmp1604;
    assign tmp1635 = tmp1633 | tmp1674;
    assign tmp1636 = tmp1621 & tmp1635;
    assign tmp1641 = tmp10 - tmp5375;
    assign tmp1645 = tmp2613 ^ tmp542;
    assign tmp1661 = tmp2787 & tmp2236;
    assign tmp1666 = tmp5375 - tmp1596;
    assign tmp1667 = {tmp1666[8]};
    assign tmp1670 = tmp1667 ^ tmp1604;
    assign tmp1671 = {tmp1596[7]};
    assign tmp1672 = ~tmp1671;
    assign tmp1673 = tmp1670 ^ tmp1672;
    assign tmp1674 = tmp5375 == tmp1596;
    assign tmp1675 = tmp1673 | tmp1674;
    assign tmp1676 = tmp1661 & tmp1675;
    assign tmp1677 = tmp1636 ? const_169_127 : tmp1596;
    assign tmp1678 = tmp1676 ? _ver_out_tmp_10 : tmp1677;
    assign tmp1692 = tmp1832 & tmp1833;
    assign tmp1694 = tmp1692 & tmp2111;
    assign tmp1715 = {tmp1731, tmp12};
    assign tmp1719 = tmp1715 + tmp649;
    assign tmp1720 = {tmp1719[8], tmp1719[7], tmp1719[6], tmp1719[5], tmp1719[4], tmp1719[3], tmp1719[2], tmp1719[1], tmp1719[0]};
    assign tmp1721 = {tmp1720[7], tmp1720[6], tmp1720[5], tmp1720[4], tmp1720[3], tmp1720[2], tmp1720[1], tmp1720[0]};
    assign tmp1731 = {tmp12[7]};
    assign tmp1746 = tmp1260 & tmp676;
    assign tmp1751 = tmp1721 - tmp5375;
    assign tmp1752 = {tmp1751[8]};
    assign tmp1753 = {tmp1721[7]};
    assign tmp1754 = ~tmp1753;
    assign tmp1755 = tmp1752 ^ tmp1754;
    assign tmp1758 = tmp1755 ^ tmp1604;
    assign tmp1759 = tmp1721 == tmp5375;
    assign tmp1760 = tmp1758 | tmp1759;
    assign tmp1761 = tmp1746 & tmp1760;
    assign tmp1766 = tmp12 - tmp5375;
    assign tmp1770 = tmp589 ^ tmp2258;
    assign tmp1778 = tmp13 - tmp5375;
    assign tmp1779 = {tmp1778[8]};
    assign tmp1781 = ~tmp711;
    assign tmp1783 = {tmp5375[7]};
    assign tmp1786 = tmp595 & tmp2274;
    assign tmp1791 = tmp5375 - tmp1721;
    assign tmp1792 = {tmp1791[8]};
    assign tmp1795 = tmp1792 ^ tmp1604;
    assign tmp1798 = tmp1795 ^ tmp1754;
    assign tmp1800 = tmp1798 | tmp1759;
    assign tmp1801 = tmp1786 & tmp1800;
    assign tmp1802 = tmp1761 ? const_177_127 : tmp1721;
    assign tmp1803 = tmp1801 ? _ver_out_tmp_58 : tmp1802;
    assign tmp1820 = tmp1694 & tmp1587;
    assign tmp1832 = tmp1545 & tmp2081;
    assign tmp1833 = ~tmp1177;
    assign tmp1844 = tmp767 + tmp888;
    assign tmp1845 = {tmp1844[8], tmp1844[7], tmp1844[6], tmp1844[5], tmp1844[4], tmp1844[3], tmp1844[2], tmp1844[1], tmp1844[0]};
    assign tmp1846 = {tmp1845[7], tmp1845[6], tmp1845[5], tmp1845[4], tmp1845[3], tmp1845[2], tmp1845[1], tmp1845[0]};
    assign tmp1858 = tmp281 ^ tmp283;
    assign tmp1870 = tmp348 ^ tmp942;
    assign tmp1871 = tmp1858 & tmp1870;
    assign tmp1876 = tmp1846 - tmp5375;
    assign tmp1877 = {tmp1876[8]};
    assign tmp1878 = {tmp1846[7]};
    assign tmp1880 = tmp1877 ^ tmp1922;
    assign tmp1883 = tmp1880 ^ tmp1604;
    assign tmp1884 = tmp1846 == tmp5375;
    assign tmp1885 = tmp1883 | tmp1884;
    assign tmp1886 = tmp1871 & tmp1885;
    assign tmp1893 = {tmp14[7]};
    assign tmp1907 = tmp7426 ^ tmp942;
    assign tmp1911 = tmp7356 & tmp2323;
    assign tmp1916 = tmp5375 - tmp1846;
    assign tmp1917 = {tmp1916[8]};
    assign tmp1920 = tmp1917 ^ tmp1604;
    assign tmp1922 = ~tmp1878;
    assign tmp1923 = tmp1920 ^ tmp1922;
    assign tmp1925 = tmp1923 | tmp1884;
    assign tmp1926 = tmp1911 & tmp1925;
    assign tmp1927 = tmp1886 ? const_185_127 : tmp1846;
    assign tmp1928 = tmp1926 ? _ver_out_tmp_14 : tmp1927;
    assign tmp1953 = tmp4780 & tmp1110;
    assign tmp1968 = {tmp7579, tmp17};
    assign tmp1969 = tmp770 + tmp1968;
    assign tmp1970 = {tmp1969[8], tmp1969[7], tmp1969[6], tmp1969[5], tmp1969[4], tmp1969[3], tmp1969[2], tmp1969[1], tmp1969[0]};
    assign tmp1971 = {tmp1970[7], tmp1970[6], tmp1970[5], tmp1970[4], tmp1970[3], tmp1970[2], tmp1970[1], tmp1970[0]};
    assign tmp1996 = tmp7483 & tmp918;
    assign tmp2001 = tmp1971 - tmp5375;
    assign tmp2002 = {tmp2001[8]};
    assign tmp2003 = {tmp1971[7]};
    assign tmp2004 = ~tmp2003;
    assign tmp2005 = tmp2002 ^ tmp2004;
    assign tmp2008 = tmp2005 ^ tmp1604;
    assign tmp2010 = tmp2008 | tmp2049;
    assign tmp2011 = tmp1996 & tmp2010;
    assign tmp2019 = ~tmp1396;
    assign tmp2036 = tmp7508 & tmp7584;
    assign tmp2041 = tmp5375 - tmp1971;
    assign tmp2042 = {tmp2041[8]};
    assign tmp2045 = tmp2042 ^ tmp1604;
    assign tmp2048 = tmp2045 ^ tmp2004;
    assign tmp2049 = tmp5375 == tmp1971;
    assign tmp2050 = tmp2048 | tmp2049;
    assign tmp2051 = tmp2036 & tmp2050;
    assign tmp2052 = tmp2011 ? const_193_127 : tmp1971;
    assign tmp2053 = tmp2051 ? _ver_out_tmp_16 : tmp2052;
    assign tmp2081 = ~tmp1122;
    assign tmp2088 = my_calculator_in_y == const_195_8;
    assign tmp2089 = tmp10 == _ver_out_tmp_17;
    assign tmp2111 = ~tmp1460;
    assign tmp2132 = ~tmp1121;
    assign tmp2167 = ~tmp1587;
    assign tmp2169 = tmp2195 & tmp2088;
    assign tmp2195 = tmp1694 & tmp2167;
    assign tmp2198 = {const_217_0, const_216_3};
    assign tmp2199 = my_calculator_ctrl == tmp2198;
    assign tmp2224 = tmp2787 == tmp2236;
    assign tmp2229 = tmp11 - tmp5375;
    assign tmp2230 = {tmp2229[8]};
    assign tmp2236 = tmp701 ^ tmp1604;
    assign tmp2249 = tmp2236 == tmp595;
    assign tmp2250 = tmp2224 & tmp2249;
    assign tmp2258 = ~tmp1731;
    assign tmp2265 = {const_223_0, const_223_0, const_223_0, const_223_0, const_223_0, const_223_0, const_223_0};
    assign tmp2274 = tmp713 ^ tmp1604;
    assign tmp2275 = tmp595 == tmp2274;
    assign tmp2276 = tmp2250 & tmp2275;
    assign tmp2311 = tmp7356 == tmp2323;
    assign tmp2323 = tmp1907 ^ tmp1604;
    assign tmp2336 = tmp2323 == tmp7508;
    assign tmp2337 = tmp2311 & tmp2336;
    assign tmp2355 = {tmp951[8]};
    assign tmp2362 = tmp7508 == tmp7584;
    assign tmp2363 = tmp2337 & tmp2362;
    assign tmp2376 = tmp14 == tmp5375;
    assign tmp2379 = tmp15 == tmp5375;
    assign tmp2380 = tmp2376 | tmp2379;
    assign tmp2384 = tmp2380 | tmp2748;
    assign tmp2387 = tmp17 == tmp5375;
    assign tmp2388 = tmp2384 | tmp2387;
    assign tmp2399 = tmp7862 & tmp7863;
    assign tmp2400 = ~tmp7864;
    assign tmp2401 = tmp2399 & tmp2400;
    assign tmp2412 = {tmp10[0]};
    assign tmp2413 = {tmp11[0]};
    assign tmp2414 = tmp2412 | tmp2413;
    assign tmp2415 = {tmp12[0]};
    assign tmp2416 = tmp2414 | tmp2415;
    assign tmp2417 = {tmp13[0]};
    assign tmp2418 = tmp2416 | tmp2417;
    assign tmp2419 = ~tmp2418;
    assign tmp2442 = tmp7865 & tmp2787;
    assign tmp2455 = tmp2442 & tmp7356;
    assign tmp2481 = tmp6763 ? tmp4109 : tmp657;
    assign tmp2482 = {tmp2481[7], tmp2481[6], tmp2481[5], tmp2481[4], tmp2481[3], tmp2481[2], tmp2481[1], tmp2481[0]};
    assign tmp2500 = tmp6798 ? tmp4109 : tmp548;
    assign tmp2501 = {tmp2500[7], tmp2500[6], tmp2500[5], tmp2500[4], tmp2500[3], tmp2500[2], tmp2500[1], tmp2500[0]};
    assign tmp2512 = tmp2549 & tmp2455;
    assign tmp2516 = tmp5375 - tmp13;
    assign tmp2520 = {tmp7157[7], tmp7157[6], tmp7157[5], tmp7157[4], tmp7157[3], tmp7157[2], tmp7157[1], tmp7157[0]};
    assign tmp2532 = tmp14 == _ver_out_tmp_29;
    assign tmp2539 = {tmp1064[7], tmp1064[6], tmp1064[5], tmp1064[4], tmp1064[3], tmp1064[2], tmp1064[1], tmp1064[0]};
    assign tmp2549 = tmp5036 & tmp2199;
    assign tmp2558 = {tmp1089[7], tmp1089[6], tmp1089[5], tmp1089[4], tmp1089[3], tmp1089[2], tmp1089[1], tmp1089[0]};
    assign tmp2573 = tmp5375 - tmp16;
    assign tmp2577 = {tmp6816[7], tmp6816[6], tmp6816[5], tmp6816[4], tmp6816[3], tmp6816[2], tmp6816[1], tmp6816[0]};
    assign tmp2585 = ~tmp1110;
    assign tmp2589 = tmp17 == _ver_out_tmp_34;
    assign tmp2595 = tmp2589 ? tmp4109 : tmp6848;
    assign tmp2596 = {tmp2595[7], tmp2595[6], tmp2595[5], tmp2595[4], tmp2595[3], tmp2595[2], tmp2595[1], tmp2595[0]};
    assign tmp2613 = {tmp1641[8]};
    assign tmp2624 = tmp14 - tmp5375;
    assign tmp2632 = tmp2787 & tmp7356;
    assign tmp2633 = ~tmp2632;
    assign tmp2634 = tmp7865 & tmp2633;
    assign tmp2659 = tmp2549 & tmp2671;
    assign tmp2660 = tmp2659 & tmp2634;
    assign tmp2671 = ~tmp2455;
    assign tmp2745 = tmp2376 & tmp2379;
    assign tmp2748 = tmp16 == tmp5375;
    assign tmp2749 = tmp2745 & tmp2748;
    assign tmp2753 = tmp2749 & tmp2387;
    assign tmp2764 = tmp2549 & tmp2753;
    assign tmp2787 = tmp1645 ^ tmp1604;
    assign tmp2800 = tmp2787 == tmp7356;
    assign tmp2801 = ~tmp2800;
    assign tmp2895 = tmp3054 & tmp2801;
    assign tmp2918 = {tmp7870[7], tmp7870[6], tmp7870[5], tmp7870[4], tmp7870[3], tmp7870[2], tmp7870[1]};
    assign tmp2919 = {tmp2918[6]};
    assign tmp2921 = {tmp2919, tmp2918};
    assign tmp2924 = tmp7886 - tmp2921;
    assign tmp2925 = {tmp2924[8]};
    assign tmp2927 = ~tmp3596;
    assign tmp2928 = tmp2925 ^ tmp2927;
    assign tmp2931 = tmp2928 ^ tmp5530;
    assign tmp2932 = tmp2921 == tmp7886;
    assign tmp2933 = tmp2931 | tmp2932;
    assign tmp2935 = {tmp4848[6]};
    assign tmp2937 = {tmp2935, tmp4848};
    assign tmp2940 = tmp7890 - tmp2937;
    assign tmp2941 = {tmp2940[8]};
    assign tmp2944 = tmp2941 ^ tmp3612;
    assign tmp2947 = tmp2944 ^ tmp5686;
    assign tmp2948 = tmp2937 == tmp7890;
    assign tmp2949 = tmp2947 | tmp2948;
    assign tmp2950 = tmp2933 & tmp2949;
    assign tmp2957 = tmp7894 - tmp3062;
    assign tmp2958 = {tmp2957[8]};
    assign tmp2959 = {tmp3062[7]};
    assign tmp2960 = ~tmp2959;
    assign tmp2961 = tmp2958 ^ tmp2960;
    assign tmp2964 = tmp2961 ^ tmp3401;
    assign tmp2965 = tmp3062 == tmp7894;
    assign tmp2966 = tmp2964 | tmp2965;
    assign tmp2967 = tmp2950 & tmp2966;
    assign tmp2968 = {tmp7882[7], tmp7882[6], tmp7882[5], tmp7882[4], tmp7882[3], tmp7882[2], tmp7882[1]};
    assign tmp2974 = tmp7898 - tmp3083;
    assign tmp2975 = {tmp2974[8]};
    assign tmp2977 = ~tmp3641;
    assign tmp2978 = tmp2975 ^ tmp2977;
    assign tmp2981 = tmp2978 ^ tmp3497;
    assign tmp2982 = tmp3083 == tmp7898;
    assign tmp2983 = tmp2981 | tmp2982;
    assign tmp2984 = tmp2967 & tmp2983;
    assign tmp3054 = tmp7385 & tmp7865;
    assign tmp3062 = {tmp4877, tmp3618};
    assign tmp3079 = tmp3150 & tmp7866;
    assign tmp3081 = {tmp2968[6]};
    assign tmp3083 = {tmp3081, tmp2968};
    assign tmp3115 = tmp3054 & tmp6025;
    assign tmp3150 = tmp3115 & tmp2984;
    assign tmp3222 = tmp3150 & tmp3387;
    assign tmp3241 = {tmp7886[6], tmp7886[5], tmp7886[4], tmp7886[3], tmp7886[2], tmp7886[1], tmp7886[0]};
    assign tmp3259 = tmp5129 - tmp5375;
    assign tmp3261 = {tmp5129[7]};
    assign tmp3279 = tmp5553 ^ tmp1604;
    assign tmp3284 = tmp5375 - tmp5129;
    assign tmp3285 = {tmp3284[8]};
    assign tmp3290 = ~tmp3261;
    assign tmp3293 = tmp5568 | tmp5569;
    assign tmp3316 = {tmp5652, const_325_0};
    assign tmp3337 = tmp5228 ^ tmp3364;
    assign tmp3364 = ~tmp5229;
    assign tmp3367 = tmp5259 | tmp5703;
    assign tmp3368 = tmp4589 & tmp3367;
    assign tmp3369 = tmp5678 ? const_330_127 : tmp3316;
    assign tmp3370 = tmp3368 ? _ver_out_tmp_60 : tmp3369;
    assign tmp3387 = ~tmp7866;
    assign tmp3395 = tmp5375 - tmp7894;
    assign tmp3399 = tmp5793 ^ tmp1604;
    assign tmp3400 = {tmp7894[7]};
    assign tmp3401 = ~tmp3400;
    assign tmp3408 = {tmp5308[8]};
    assign tmp3411 = tmp3408 ^ tmp5835;
    assign tmp3415 = tmp4642 & tmp5315;
    assign tmp3424 = tmp5322 ^ tmp3401;
    assign tmp3427 = tmp3424 ^ tmp1604;
    assign tmp3432 = tmp5375 - tmp5291;
    assign tmp3436 = tmp5334 ^ tmp1604;
    assign tmp3439 = tmp3436 ^ tmp5835;
    assign tmp3444 = tmp5343 ? _ver_out_tmp_62 : tmp5840;
    assign tmp3470 = {tmp5377[8]};
    assign tmp3489 = tmp5384 & tmp5945;
    assign tmp3494 = tmp7898 - tmp5375;
    assign tmp3497 = ~tmp5404;
    assign tmp3512 = ~tmp5391;
    assign tmp3513 = tmp5418 ^ tmp3512;
    assign tmp3514 = tmp5375 == tmp5372;
    assign tmp3518 = tmp5424 ? _ver_out_tmp_66 : tmp5425;
    assign tmp3543 = tmp4466 ^ tmp3728;
    assign tmp3544 = {tmp7886[7]};
    assign tmp3546 = tmp3543 ^ tmp5530;
    assign tmp3547 = tmp7870 == tmp7886;
    assign tmp3548 = tmp3546 | tmp3547;
    assign tmp3552 = {tmp4542[8]};
    assign tmp3555 = tmp3552 ^ tmp5713;
    assign tmp3558 = tmp3555 ^ tmp5686;
    assign tmp3559 = tmp7874 == tmp7890;
    assign tmp3560 = tmp3558 | tmp3559;
    assign tmp3561 = tmp3548 & tmp3560;
    assign tmp3566 = {tmp7878[7]};
    assign tmp3567 = ~tmp3566;
    assign tmp3568 = tmp4621 ^ tmp3567;
    assign tmp3571 = tmp3568 ^ tmp3401;
    assign tmp3572 = tmp7878 == tmp7894;
    assign tmp3573 = tmp3571 | tmp3572;
    assign tmp3574 = tmp3561 & tmp3573;
    assign tmp3577 = tmp7898 - tmp7882;
    assign tmp3581 = tmp4699 ^ tmp5887;
    assign tmp3584 = tmp3581 ^ tmp3497;
    assign tmp3585 = tmp7882 == tmp7898;
    assign tmp3586 = tmp3584 | tmp3585;
    assign tmp3587 = tmp3574 & tmp3586;
    assign tmp3594 = tmp2921 - tmp7886;
    assign tmp3595 = {tmp3594[8]};
    assign tmp3596 = {tmp2921[7]};
    assign tmp3598 = tmp3595 ^ tmp2927;
    assign tmp3601 = tmp3598 ^ tmp5530;
    assign tmp3602 = tmp3587 & tmp3601;
    assign tmp3609 = tmp2937 - tmp7890;
    assign tmp3610 = {tmp3609[8]};
    assign tmp3611 = {tmp2937[7]};
    assign tmp3612 = ~tmp3611;
    assign tmp3613 = tmp3610 ^ tmp3612;
    assign tmp3616 = tmp3613 ^ tmp5686;
    assign tmp3617 = tmp3602 & tmp3616;
    assign tmp3618 = {tmp7878[7], tmp7878[6], tmp7878[5], tmp7878[4], tmp7878[3], tmp7878[2], tmp7878[1]};
    assign tmp3624 = tmp3062 - tmp7894;
    assign tmp3625 = {tmp3624[8]};
    assign tmp3628 = tmp3625 ^ tmp2960;
    assign tmp3631 = tmp3628 ^ tmp3401;
    assign tmp3632 = tmp3617 & tmp3631;
    assign tmp3639 = tmp3083 - tmp7898;
    assign tmp3640 = {tmp3639[8]};
    assign tmp3641 = {tmp3083[7]};
    assign tmp3643 = tmp3640 ^ tmp2977;
    assign tmp3646 = tmp3643 ^ tmp3497;
    assign tmp3647 = tmp3632 & tmp3646;
    assign tmp3701 = tmp4218 & tmp3647;
    assign tmp3702 = _ver_out_tmp_68 == tmp7886;
    assign tmp3708 = tmp3702 ? tmp4109 : tmp5134;
    assign tmp3711 = {tmp6070, tmp7870};
    assign tmp3712 = {tmp3708[8]};
    assign tmp3722 = tmp5375 - tmp7870;
    assign tmp3728 = ~tmp3764;
    assign tmp3735 = {tmp6094[9]};
    assign tmp3740 = ~tmp3712;
    assign tmp3741 = tmp6098 ^ tmp3740;
    assign tmp3742 = tmp6089 & tmp3741;
    assign tmp3747 = tmp6077 - tmp5375;
    assign tmp3749 = {tmp6077[7]};
    assign tmp3751 = tmp6108 ^ tmp6153;
    assign tmp3754 = tmp3751 ^ tmp1604;
    assign tmp3757 = tmp3742 & tmp6116;
    assign tmp3764 = {tmp7870[7]};
    assign tmp3778 = tmp6135 ^ tmp3740;
    assign tmp3788 = {tmp6147[8]};
    assign tmp3794 = tmp6151 ^ tmp6153;
    assign tmp3795 = tmp5375 == tmp6077;
    assign tmp3796 = tmp3794 | tmp3795;
    assign tmp3797 = tmp6142 & tmp3796;
    assign tmp3799 = tmp3797 ? _ver_out_tmp_75 : tmp6158;
    assign tmp3842 = tmp6210 ? tmp4109 : tmp5215;
    assign tmp3844 = {tmp4547, tmp4547};
    assign tmp3846 = {tmp3842[8]};
    assign tmp3856 = tmp5375 - tmp7874;
    assign tmp3857 = {tmp3856[8]};
    assign tmp3860 = tmp3857 ^ tmp1604;
    assign tmp3874 = ~tmp3846;
    assign tmp3875 = tmp6246 ^ tmp3874;
    assign tmp3876 = tmp5598 & tmp3875;
    assign tmp3885 = tmp6256 ^ tmp3927;
    assign tmp3888 = tmp3885 ^ tmp1604;
    assign tmp3890 = tmp3888 | tmp6303;
    assign tmp3891 = tmp3876 & tmp3890;
    assign tmp3908 = tmp3842 - tmp4041;
    assign tmp3912 = tmp6283 ^ tmp3874;
    assign tmp3913 = {tmp4041[8]};
    assign tmp3915 = tmp3912 ^ tmp6140;
    assign tmp3916 = tmp6277 & tmp3915;
    assign tmp3922 = {tmp6295[8]};
    assign tmp3925 = tmp3922 ^ tmp1604;
    assign tmp3926 = {tmp6225[7]};
    assign tmp3927 = ~tmp3926;
    assign tmp3931 = tmp3916 & tmp6304;
    assign tmp3933 = tmp3931 ? _ver_out_tmp_85 : tmp6306;
    assign tmp3976 = tmp6358 ? tmp4109 : tmp3395;
    assign tmp3991 = {tmp5725[8]};
    assign tmp3994 = tmp3991 ^ tmp1604;
    assign tmp4002 = tmp4041 - tmp3976;
    assign tmp4006 = tmp6391 ^ tmp6140;
    assign tmp4007 = {tmp3976[8]};
    assign tmp4015 = tmp6373 - tmp5375;
    assign tmp4016 = {tmp4015[8]};
    assign tmp4019 = tmp4016 ^ tmp4061;
    assign tmp4022 = tmp4019 ^ tmp1604;
    assign tmp4024 = tmp4022 | tmp4063;
    assign tmp4025 = tmp6398 & tmp4024;
    assign tmp4037 = tmp5754 ^ tmp1604;
    assign tmp4041 = {tmp6387, const_383_0};
    assign tmp4042 = tmp3976 - tmp4041;
    assign tmp4045 = ~tmp4007;
    assign tmp4046 = tmp6431 ^ tmp4045;
    assign tmp4050 = tmp4037 & tmp6437;
    assign tmp4056 = {tmp6443[8]};
    assign tmp4059 = tmp4056 ^ tmp1604;
    assign tmp4061 = ~tmp6405;
    assign tmp4062 = tmp4059 ^ tmp4061;
    assign tmp4063 = tmp5375 == tmp6373;
    assign tmp4064 = tmp4062 | tmp4063;
    assign tmp4065 = tmp4050 & tmp4064;
    assign tmp4067 = tmp4065 ? _ver_out_tmp_27 : tmp6454;
    assign tmp4109 = {tmp133, const_390_127};
    assign tmp4110 = tmp6506 ? tmp4109 : tmp5377;
    assign tmp4116 = {tmp6516, tmp4110};
    assign tmp4118 = {tmp6519[9], tmp6519[8], tmp6519[7], tmp6519[6], tmp6519[5], tmp6519[4], tmp6519[3], tmp6519[2], tmp6519[1], tmp6519[0]};
    assign tmp4119 = {tmp4118[7], tmp4118[6], tmp4118[5], tmp4118[4], tmp4118[3], tmp4118[2], tmp4118[1], tmp4118[0]};
    assign tmp4125 = {tmp5859[8]};
    assign tmp4128 = tmp4125 ^ tmp1604;
    assign tmp4136 = tmp4041 - tmp4110;
    assign tmp4143 = tmp6542 ^ tmp6544;
    assign tmp4144 = tmp6533 & tmp4143;
    assign tmp4156 = tmp6555 ^ tmp1604;
    assign tmp4157 = tmp4119 == tmp5375;
    assign tmp4158 = tmp4156 | tmp4157;
    assign tmp4159 = tmp4144 & tmp4158;
    assign tmp4176 = tmp4110 - tmp4041;
    assign tmp4180 = tmp6579 ^ tmp6544;
    assign tmp4183 = tmp4180 ^ tmp6140;
    assign tmp4184 = tmp6573 & tmp4183;
    assign tmp4189 = tmp5375 - tmp4119;
    assign tmp4190 = {tmp4189[8]};
    assign tmp4193 = tmp4190 ^ tmp1604;
    assign tmp4194 = {tmp4119[7]};
    assign tmp4196 = tmp4193 ^ tmp6597;
    assign tmp4198 = tmp4196 | tmp4157;
    assign tmp4200 = tmp4159 ? const_398_127 : tmp4119;
    assign tmp4201 = tmp6601 ? _ver_out_tmp_33 : tmp4200;
    assign tmp4218 = tmp3115 & tmp4358;
    assign tmp4222 = tmp7870 - tmp7886;
    assign tmp4223 = {tmp4222[8]};
    assign tmp4226 = tmp4223 ^ tmp3728;
    assign tmp4229 = tmp4226 ^ tmp5530;
    assign tmp4232 = tmp7874 - tmp7890;
    assign tmp4233 = {tmp4232[8]};
    assign tmp4236 = tmp4233 ^ tmp5713;
    assign tmp4239 = tmp4236 ^ tmp5686;
    assign tmp4240 = tmp4229 & tmp4239;
    assign tmp4243 = tmp7878 - tmp7894;
    assign tmp4244 = {tmp4243[8]};
    assign tmp4247 = tmp4244 ^ tmp3567;
    assign tmp4250 = tmp4247 ^ tmp3401;
    assign tmp4251 = tmp4240 & tmp4250;
    assign tmp4254 = tmp7882 - tmp7898;
    assign tmp4255 = {tmp4254[8]};
    assign tmp4258 = tmp4255 ^ tmp5887;
    assign tmp4261 = tmp4258 ^ tmp3497;
    assign tmp4262 = tmp4251 & tmp4261;
    assign tmp4280 = ~tmp3647;
    assign tmp4358 = ~tmp2984;
    assign tmp4362 = tmp6030 & tmp4262;
    assign tmp4465 = tmp7886 - tmp7870;
    assign tmp4466 = {tmp4465[8]};
    assign tmp4469 = tmp4466 ^ tmp5530;
    assign tmp4472 = tmp4469 ^ tmp3728;
    assign tmp4473 = {tmp7886[5], tmp7886[4], tmp7886[3], tmp7886[2], tmp7886[1], tmp7886[0]};
    assign tmp4474 = {tmp4473, const_402_0};
    assign tmp4483 = tmp5135 ^ tmp1604;
    assign tmp4486 = tmp4483 ^ tmp5530;
    assign tmp4491 = tmp4474 - tmp5375;
    assign tmp4492 = {tmp4491[8]};
    assign tmp4495 = tmp4492 ^ tmp4522;
    assign tmp4498 = tmp4495 ^ tmp1604;
    assign tmp4499 = tmp4486 & tmp4498;
    assign tmp4505 = {tmp5549[8]};
    assign tmp4516 = tmp5375 - tmp4474;
    assign tmp4517 = {tmp4516[8]};
    assign tmp4520 = tmp4517 ^ tmp1604;
    assign tmp4521 = {tmp4474[7]};
    assign tmp4522 = ~tmp4521;
    assign tmp4523 = tmp4520 ^ tmp4522;
    assign tmp4524 = tmp5375 == tmp4474;
    assign tmp4525 = tmp4523 | tmp4524;
    assign tmp4526 = tmp3279 & tmp4525;
    assign tmp4527 = tmp4499 ? const_407_127 : tmp4474;
    assign tmp4528 = tmp4526 ? _ver_out_tmp_37 : tmp4527;
    assign tmp4531 = tmp7870 - tmp4528;
    assign tmp4532 = {tmp4531[8]};
    assign tmp4535 = tmp4532 ^ tmp3728;
    assign tmp4536 = {tmp4528[7]};
    assign tmp4537 = ~tmp4536;
    assign tmp4538 = tmp4535 ^ tmp4537;
    assign tmp4539 = tmp4472 & tmp4538;
    assign tmp4542 = tmp7890 - tmp7874;
    assign tmp4546 = tmp3552 ^ tmp5686;
    assign tmp4547 = {tmp7874[7]};
    assign tmp4549 = tmp4546 ^ tmp5713;
    assign tmp4550 = tmp4539 & tmp4549;
    assign tmp4551 = {tmp7890[5], tmp7890[4], tmp7890[3], tmp7890[2], tmp7890[1], tmp7890[0]};
    assign tmp4552 = {tmp4551, const_409_0};
    assign tmp4558 = {tmp5215[8]};
    assign tmp4561 = tmp4558 ^ tmp1604;
    assign tmp4564 = tmp4561 ^ tmp5686;
    assign tmp4569 = tmp4552 - tmp5375;
    assign tmp4570 = {tmp4569[8]};
    assign tmp4571 = {tmp4552[7]};
    assign tmp4572 = ~tmp4571;
    assign tmp4573 = tmp4570 ^ tmp4572;
    assign tmp4576 = tmp4573 ^ tmp1604;
    assign tmp4577 = tmp4564 & tmp4576;
    assign tmp4589 = tmp5244 ^ tmp1604;
    assign tmp4594 = tmp5375 - tmp4552;
    assign tmp4595 = {tmp4594[8]};
    assign tmp4598 = tmp4595 ^ tmp1604;
    assign tmp4601 = tmp4598 ^ tmp4572;
    assign tmp4602 = tmp5375 == tmp4552;
    assign tmp4603 = tmp4601 | tmp4602;
    assign tmp4604 = tmp4589 & tmp4603;
    assign tmp4605 = tmp4577 ? const_414_127 : tmp4552;
    assign tmp4606 = tmp4604 ? _ver_out_tmp_38 : tmp4605;
    assign tmp4609 = tmp7874 - tmp4606;
    assign tmp4610 = {tmp4609[8]};
    assign tmp4613 = tmp4610 ^ tmp5713;
    assign tmp4614 = {tmp4606[7]};
    assign tmp4615 = ~tmp4614;
    assign tmp4616 = tmp4613 ^ tmp4615;
    assign tmp4617 = tmp4550 & tmp4616;
    assign tmp4620 = tmp7894 - tmp7878;
    assign tmp4621 = {tmp4620[8]};
    assign tmp4624 = tmp4621 ^ tmp3401;
    assign tmp4627 = tmp4624 ^ tmp3567;
    assign tmp4628 = tmp4617 & tmp4627;
    assign tmp4629 = {tmp7894[5], tmp7894[4], tmp7894[3], tmp7894[2], tmp7894[1], tmp7894[0]};
    assign tmp4630 = {tmp4629, const_416_0};
    assign tmp4642 = tmp3399 ^ tmp3401;
    assign tmp4647 = tmp4630 - tmp5375;
    assign tmp4648 = {tmp4647[8]};
    assign tmp4651 = tmp4648 ^ tmp4678;
    assign tmp4654 = tmp4651 ^ tmp1604;
    assign tmp4655 = tmp4642 & tmp4654;
    assign tmp4660 = tmp7894 - tmp5375;
    assign tmp4672 = tmp5375 - tmp4630;
    assign tmp4673 = {tmp4672[8]};
    assign tmp4676 = tmp4673 ^ tmp1604;
    assign tmp4677 = {tmp4630[7]};
    assign tmp4678 = ~tmp4677;
    assign tmp4679 = tmp4676 ^ tmp4678;
    assign tmp4680 = tmp5375 == tmp4630;
    assign tmp4681 = tmp4679 | tmp4680;
    assign tmp4682 = tmp3427 & tmp4681;
    assign tmp4683 = tmp4655 ? const_421_127 : tmp4630;
    assign tmp4684 = tmp4682 ? _ver_out_tmp_41 : tmp4683;
    assign tmp4687 = tmp7878 - tmp4684;
    assign tmp4688 = {tmp4687[8]};
    assign tmp4691 = tmp4688 ^ tmp3567;
    assign tmp4692 = {tmp4684[7]};
    assign tmp4693 = ~tmp4692;
    assign tmp4694 = tmp4691 ^ tmp4693;
    assign tmp4695 = tmp4628 & tmp4694;
    assign tmp4699 = {tmp3577[8]};
    assign tmp4702 = tmp4699 ^ tmp3497;
    assign tmp4703 = {tmp7882[7]};
    assign tmp4705 = tmp4702 ^ tmp5887;
    assign tmp4706 = tmp4695 & tmp4705;
    assign tmp4707 = {tmp7898[5], tmp7898[4], tmp7898[3], tmp7898[2], tmp7898[1], tmp7898[0]};
    assign tmp4708 = {tmp4707, const_423_0};
    assign tmp4717 = tmp3470 ^ tmp1604;
    assign tmp4725 = tmp4708 - tmp5375;
    assign tmp4726 = {tmp4725[8]};
    assign tmp4727 = {tmp4708[7]};
    assign tmp4729 = tmp4726 ^ tmp4756;
    assign tmp4732 = tmp4729 ^ tmp1604;
    assign tmp4733 = tmp5384 & tmp4732;
    assign tmp4745 = tmp5406 ^ tmp1604;
    assign tmp4750 = tmp5375 - tmp4708;
    assign tmp4751 = {tmp4750[8]};
    assign tmp4754 = tmp4751 ^ tmp1604;
    assign tmp4756 = ~tmp4727;
    assign tmp4757 = tmp4754 ^ tmp4756;
    assign tmp4758 = tmp5375 == tmp4708;
    assign tmp4759 = tmp4757 | tmp4758;
    assign tmp4760 = tmp4745 & tmp4759;
    assign tmp4761 = tmp4733 ? const_428_127 : tmp4708;
    assign tmp4762 = tmp4760 ? _ver_out_tmp_43 : tmp4761;
    assign tmp4765 = tmp7882 - tmp4762;
    assign tmp4766 = {tmp4765[8]};
    assign tmp4769 = tmp4766 ^ tmp5887;
    assign tmp4770 = {tmp4762[7]};
    assign tmp4771 = ~tmp4770;
    assign tmp4772 = tmp4769 ^ tmp4771;
    assign tmp4773 = tmp4706 & tmp4772;
    assign tmp4780 = tmp1070 & tmp6951;
    assign tmp4796 = tmp6353 & tmp4773;
    assign tmp4798 = ~tmp35;
    assign tmp4848 = {tmp7874[7], tmp7874[6], tmp7874[5], tmp7874[4], tmp7874[3], tmp7874[2], tmp7874[1]};
    assign tmp4877 = {tmp3618[6]};
    assign tmp4931 = tmp4796 & tmp7866;
    assign tmp5036 = tmp4780 & tmp2585;
    assign tmp5077 = tmp4796 & tmp3387;
    assign tmp5081 = ~tmp36;
    assign tmp5129 = {tmp3241, const_432_0};
    assign tmp5134 = tmp5375 - tmp7886;
    assign tmp5135 = {tmp5134[8]};
    assign tmp5150 = tmp5537 ^ tmp3290;
    assign tmp5154 = tmp4486 & tmp5543;
    assign tmp5175 = tmp3285 ^ tmp1604;
    assign tmp5182 = tmp5154 ? const_437_127 : tmp5129;
    assign tmp5183 = tmp5571 ? _ver_out_tmp_47 : tmp5182;
    assign tmp5215 = tmp5375 - tmp7890;
    assign tmp5227 = tmp3316 - tmp5375;
    assign tmp5228 = {tmp5227[8]};
    assign tmp5229 = {tmp3316[7]};
    assign tmp5241 = {tmp5683[8]};
    assign tmp5244 = tmp5241 ^ tmp5686;
    assign tmp5253 = {tmp5695[8]};
    assign tmp5256 = tmp5253 ^ tmp1604;
    assign tmp5259 = tmp5256 ^ tmp3364;
    assign tmp5290 = {tmp7894[6], tmp7894[5], tmp7894[4], tmp7894[3], tmp7894[2], tmp7894[1], tmp7894[0]};
    assign tmp5291 = {tmp5290, const_446_0};
    assign tmp5308 = tmp5291 - tmp5375;
    assign tmp5310 = {tmp5291[7]};
    assign tmp5315 = tmp3411 ^ tmp1604;
    assign tmp5322 = {tmp4660[8]};
    assign tmp5334 = {tmp3432[8]};
    assign tmp5341 = tmp5375 == tmp5291;
    assign tmp5342 = tmp3439 | tmp5341;
    assign tmp5343 = tmp3427 & tmp5342;
    assign tmp5372 = {tmp5920, const_453_0};
    assign tmp5375 = {tmp2265, const_454_0};
    assign tmp5377 = tmp5375 - tmp7898;
    assign tmp5384 = tmp4717 ^ tmp3497;
    assign tmp5390 = {tmp5938[8]};
    assign tmp5391 = {tmp5372[7]};
    assign tmp5404 = {tmp7898[7]};
    assign tmp5406 = tmp5952 ^ tmp3497;
    assign tmp5418 = tmp5964 ^ tmp1604;
    assign tmp5424 = tmp4745 & tmp5972;
    assign tmp5425 = tmp3489 ? const_458_127 : tmp5372;
    assign tmp5452 = {tmp7870[6], tmp7870[5], tmp7870[4], tmp7870[3], tmp7870[2], tmp7870[1], tmp7870[0]};
    assign tmp5453 = {tmp5452, const_460_0};
    assign tmp5459 = {tmp3722[8]};
    assign tmp5470 = tmp5453 - tmp5375;
    assign tmp5471 = {tmp5470[8]};
    assign tmp5473 = ~tmp5500;
    assign tmp5474 = tmp5471 ^ tmp5473;
    assign tmp5477 = tmp5474 ^ tmp1604;
    assign tmp5478 = tmp6089 & tmp5477;
    assign tmp5483 = tmp7870 - tmp5375;
    assign tmp5495 = tmp5375 - tmp5453;
    assign tmp5496 = {tmp5495[8]};
    assign tmp5499 = tmp5496 ^ tmp1604;
    assign tmp5500 = {tmp5453[7]};
    assign tmp5502 = tmp5499 ^ tmp5473;
    assign tmp5503 = tmp5375 == tmp5453;
    assign tmp5504 = tmp5502 | tmp5503;
    assign tmp5505 = tmp6129 & tmp5504;
    assign tmp5506 = tmp5478 ? const_465_127 : tmp5453;
    assign tmp5507 = tmp5505 ? _ver_out_tmp_90 : tmp5506;
    assign tmp5510 = tmp7886 - tmp5507;
    assign tmp5511 = {tmp5510[8]};
    assign tmp5514 = tmp5511 ^ tmp5530;
    assign tmp5515 = {tmp5507[7]};
    assign tmp5516 = ~tmp5515;
    assign tmp5517 = tmp5514 ^ tmp5516;
    assign tmp5530 = ~tmp3544;
    assign tmp5537 = {tmp3259[8]};
    assign tmp5543 = tmp5150 ^ tmp1604;
    assign tmp5549 = tmp7886 - tmp5375;
    assign tmp5553 = tmp4505 ^ tmp5530;
    assign tmp5568 = tmp5175 ^ tmp3290;
    assign tmp5569 = tmp5375 == tmp5129;
    assign tmp5571 = tmp3279 & tmp3293;
    assign tmp5576 = tmp7870 - tmp5183;
    assign tmp5577 = {tmp5576[8]};
    assign tmp5580 = tmp5577 ^ tmp3728;
    assign tmp5581 = {tmp5183[7]};
    assign tmp5582 = ~tmp5581;
    assign tmp5583 = tmp5580 ^ tmp5582;
    assign tmp5584 = tmp5517 & tmp5583;
    assign tmp5585 = {tmp7874[6], tmp7874[5], tmp7874[4], tmp7874[3], tmp7874[2], tmp7874[1], tmp7874[0]};
    assign tmp5586 = {tmp5585, const_474_0};
    assign tmp5598 = tmp3860 ^ tmp5713;
    assign tmp5603 = tmp5586 - tmp5375;
    assign tmp5604 = {tmp5603[8]};
    assign tmp5607 = tmp5604 ^ tmp5634;
    assign tmp5610 = tmp5607 ^ tmp1604;
    assign tmp5611 = tmp5598 & tmp5610;
    assign tmp5620 = tmp6271 ^ tmp5713;
    assign tmp5628 = tmp5375 - tmp5586;
    assign tmp5629 = {tmp5628[8]};
    assign tmp5632 = tmp5629 ^ tmp1604;
    assign tmp5633 = {tmp5586[7]};
    assign tmp5634 = ~tmp5633;
    assign tmp5635 = tmp5632 ^ tmp5634;
    assign tmp5636 = tmp5375 == tmp5586;
    assign tmp5637 = tmp5635 | tmp5636;
    assign tmp5638 = tmp6277 & tmp5637;
    assign tmp5639 = tmp5611 ? const_479_127 : tmp5586;
    assign tmp5640 = tmp5638 ? _ver_out_tmp_67 : tmp5639;
    assign tmp5643 = tmp7890 - tmp5640;
    assign tmp5644 = {tmp5643[8]};
    assign tmp5647 = tmp5644 ^ tmp5686;
    assign tmp5648 = {tmp5640[7]};
    assign tmp5649 = ~tmp5648;
    assign tmp5650 = tmp5647 ^ tmp5649;
    assign tmp5651 = tmp5584 & tmp5650;
    assign tmp5652 = {tmp7890[6], tmp7890[5], tmp7890[4], tmp7890[3], tmp7890[2], tmp7890[1], tmp7890[0]};
    assign tmp5677 = tmp3337 ^ tmp1604;
    assign tmp5678 = tmp4564 & tmp5677;
    assign tmp5683 = tmp7890 - tmp5375;
    assign tmp5685 = {tmp7890[7]};
    assign tmp5686 = ~tmp5685;
    assign tmp5695 = tmp5375 - tmp3316;
    assign tmp5703 = tmp5375 == tmp3316;
    assign tmp5710 = tmp7874 - tmp3370;
    assign tmp5711 = {tmp5710[8]};
    assign tmp5713 = ~tmp4547;
    assign tmp5714 = tmp5711 ^ tmp5713;
    assign tmp5715 = {tmp3370[7]};
    assign tmp5716 = ~tmp5715;
    assign tmp5717 = tmp5714 ^ tmp5716;
    assign tmp5718 = tmp5651 & tmp5717;
    assign tmp5719 = {tmp7878[6], tmp7878[5], tmp7878[4], tmp7878[3], tmp7878[2], tmp7878[1], tmp7878[0]};
    assign tmp5720 = {tmp5719, const_488_0};
    assign tmp5725 = tmp5375 - tmp7878;
    assign tmp5737 = tmp5720 - tmp5375;
    assign tmp5738 = {tmp5737[8]};
    assign tmp5741 = tmp5738 ^ tmp5768;
    assign tmp5744 = tmp5741 ^ tmp1604;
    assign tmp5745 = tmp6385 & tmp5744;
    assign tmp5750 = tmp7878 - tmp5375;
    assign tmp5754 = tmp6419 ^ tmp3567;
    assign tmp5762 = tmp5375 - tmp5720;
    assign tmp5763 = {tmp5762[8]};
    assign tmp5766 = tmp5763 ^ tmp1604;
    assign tmp5767 = {tmp5720[7]};
    assign tmp5768 = ~tmp5767;
    assign tmp5769 = tmp5766 ^ tmp5768;
    assign tmp5770 = tmp5375 == tmp5720;
    assign tmp5771 = tmp5769 | tmp5770;
    assign tmp5772 = tmp4037 & tmp5771;
    assign tmp5773 = tmp5745 ? const_493_127 : tmp5720;
    assign tmp5774 = tmp5772 ? _ver_out_tmp_74 : tmp5773;
    assign tmp5777 = tmp7894 - tmp5774;
    assign tmp5778 = {tmp5777[8]};
    assign tmp5781 = tmp5778 ^ tmp3401;
    assign tmp5782 = {tmp5774[7]};
    assign tmp5783 = ~tmp5782;
    assign tmp5784 = tmp5781 ^ tmp5783;
    assign tmp5785 = tmp5718 & tmp5784;
    assign tmp5793 = {tmp3395[8]};
    assign tmp5835 = ~tmp5310;
    assign tmp5840 = tmp3415 ? const_500_127 : tmp5291;
    assign tmp5844 = tmp7878 - tmp3444;
    assign tmp5845 = {tmp5844[8]};
    assign tmp5848 = tmp5845 ^ tmp3567;
    assign tmp5849 = {tmp3444[7]};
    assign tmp5850 = ~tmp5849;
    assign tmp5851 = tmp5848 ^ tmp5850;
    assign tmp5852 = tmp5785 & tmp5851;
    assign tmp5853 = {tmp7882[6], tmp7882[5], tmp7882[4], tmp7882[3], tmp7882[2], tmp7882[1], tmp7882[0]};
    assign tmp5854 = {tmp5853, const_502_0};
    assign tmp5859 = tmp5375 - tmp7882;
    assign tmp5871 = tmp5854 - tmp5375;
    assign tmp5872 = {tmp5871[8]};
    assign tmp5873 = {tmp5854[7]};
    assign tmp5875 = tmp5872 ^ tmp5902;
    assign tmp5878 = tmp5875 ^ tmp1604;
    assign tmp5879 = tmp6533 & tmp5878;
    assign tmp5887 = ~tmp4703;
    assign tmp5888 = tmp6567 ^ tmp5887;
    assign tmp5896 = tmp5375 - tmp5854;
    assign tmp5897 = {tmp5896[8]};
    assign tmp5900 = tmp5897 ^ tmp1604;
    assign tmp5902 = ~tmp5873;
    assign tmp5903 = tmp5900 ^ tmp5902;
    assign tmp5904 = tmp5375 == tmp5854;
    assign tmp5905 = tmp5903 | tmp5904;
    assign tmp5906 = tmp6573 & tmp5905;
    assign tmp5907 = tmp5879 ? const_507_127 : tmp5854;
    assign tmp5908 = tmp5906 ? _ver_out_tmp_82 : tmp5907;
    assign tmp5911 = tmp7898 - tmp5908;
    assign tmp5912 = {tmp5911[8]};
    assign tmp5915 = tmp5912 ^ tmp3497;
    assign tmp5916 = {tmp5908[7]};
    assign tmp5917 = ~tmp5916;
    assign tmp5918 = tmp5915 ^ tmp5917;
    assign tmp5919 = tmp5852 & tmp5918;
    assign tmp5920 = {tmp7898[6], tmp7898[5], tmp7898[4], tmp7898[3], tmp7898[2], tmp7898[1], tmp7898[0]};
    assign tmp5938 = tmp5372 - tmp5375;
    assign tmp5942 = tmp5390 ^ tmp3512;
    assign tmp5945 = tmp5942 ^ tmp1604;
    assign tmp5952 = {tmp3494[8]};
    assign tmp5963 = tmp5375 - tmp5372;
    assign tmp5964 = {tmp5963[8]};
    assign tmp5972 = tmp3513 | tmp3514;
    assign tmp5978 = tmp7882 - tmp3518;
    assign tmp5979 = {tmp5978[8]};
    assign tmp5982 = tmp5979 ^ tmp5887;
    assign tmp5983 = {tmp3518[7]};
    assign tmp5984 = ~tmp5983;
    assign tmp5985 = tmp5982 ^ tmp5984;
    assign tmp5986 = tmp5919 & tmp5985;
    assign tmp6009 = ~tmp4773;
    assign tmp6025 = ~tmp2801;
    assign tmp6030 = tmp4218 & tmp4280;
    assign tmp6070 = {tmp3764, tmp3764};
    assign tmp6074 = {tmp3712, tmp3708};
    assign tmp6075 = tmp3711 + tmp6074;
    assign tmp6076 = {tmp6075[9], tmp6075[8], tmp6075[7], tmp6075[6], tmp6075[5], tmp6075[4], tmp6075[3], tmp6075[2], tmp6075[1], tmp6075[0]};
    assign tmp6077 = {tmp6076[7], tmp6076[6], tmp6076[5], tmp6076[4], tmp6076[3], tmp6076[2], tmp6076[1], tmp6076[0]};
    assign tmp6086 = tmp5459 ^ tmp1604;
    assign tmp6089 = tmp6086 ^ tmp3728;
    assign tmp6094 = tmp4041 - tmp3708;
    assign tmp6098 = tmp3735 ^ tmp6140;
    assign tmp6108 = {tmp3747[8]};
    assign tmp6116 = tmp3754 | tmp3795;
    assign tmp6123 = {tmp5483[8]};
    assign tmp6126 = tmp6123 ^ tmp3728;
    assign tmp6129 = tmp6126 ^ tmp1604;
    assign tmp6134 = tmp3708 - tmp4041;
    assign tmp6135 = {tmp6134[9]};
    assign tmp6140 = ~tmp3913;
    assign tmp6141 = tmp3778 ^ tmp6140;
    assign tmp6142 = tmp6129 & tmp6141;
    assign tmp6147 = tmp5375 - tmp6077;
    assign tmp6151 = tmp3788 ^ tmp1604;
    assign tmp6153 = ~tmp3749;
    assign tmp6158 = tmp3757 ? const_529_127 : tmp6077;
    assign tmp6209 = tmp6356 & tmp5986;
    assign tmp6210 = _ver_out_tmp_30 == tmp7890;
    assign tmp6219 = {tmp3844, tmp7874};
    assign tmp6222 = {tmp3846, tmp3842};
    assign tmp6223 = tmp6219 + tmp6222;
    assign tmp6224 = {tmp6223[9], tmp6223[8], tmp6223[7], tmp6223[6], tmp6223[5], tmp6223[4], tmp6223[3], tmp6223[2], tmp6223[1], tmp6223[0]};
    assign tmp6225 = {tmp6224[7], tmp6224[6], tmp6224[5], tmp6224[4], tmp6224[3], tmp6224[2], tmp6224[1], tmp6224[0]};
    assign tmp6242 = tmp4041 - tmp3842;
    assign tmp6243 = {tmp6242[9]};
    assign tmp6246 = tmp6243 ^ tmp6140;
    assign tmp6255 = tmp6225 - tmp5375;
    assign tmp6256 = {tmp6255[8]};
    assign tmp6270 = tmp7874 - tmp5375;
    assign tmp6271 = {tmp6270[8]};
    assign tmp6277 = tmp5620 ^ tmp1604;
    assign tmp6283 = {tmp3908[9]};
    assign tmp6295 = tmp5375 - tmp6225;
    assign tmp6302 = tmp3925 ^ tmp3927;
    assign tmp6303 = tmp5375 == tmp6225;
    assign tmp6304 = tmp6302 | tmp6303;
    assign tmp6306 = tmp3891 ? const_542_127 : tmp6225;
    assign tmp6327 = ~tmp4262;
    assign tmp6353 = tmp6030 & tmp6327;
    assign tmp6356 = tmp6353 & tmp6009;
    assign tmp6358 = _ver_out_tmp_36 == tmp7894;
    assign tmp6366 = {tmp3566, tmp3566};
    assign tmp6367 = {tmp6366, tmp7878};
    assign tmp6370 = {tmp4007, tmp3976};
    assign tmp6371 = tmp6367 + tmp6370;
    assign tmp6372 = {tmp6371[9], tmp6371[8], tmp6371[7], tmp6371[6], tmp6371[5], tmp6371[4], tmp6371[3], tmp6371[2], tmp6371[1], tmp6371[0]};
    assign tmp6373 = {tmp6372[7], tmp6372[6], tmp6372[5], tmp6372[4], tmp6372[3], tmp6372[2], tmp6372[1], tmp6372[0]};
    assign tmp6385 = tmp3994 ^ tmp3567;
    assign tmp6387 = {const_550_0, const_550_0, const_550_0, const_550_0, const_550_0, const_550_0, const_550_0, const_550_0};
    assign tmp6391 = {tmp4002[9]};
    assign tmp6397 = tmp4006 ^ tmp4045;
    assign tmp6398 = tmp6385 & tmp6397;
    assign tmp6405 = {tmp6373[7]};
    assign tmp6419 = {tmp5750[8]};
    assign tmp6431 = {tmp4042[9]};
    assign tmp6437 = tmp4046 ^ tmp6140;
    assign tmp6443 = tmp5375 - tmp6373;
    assign tmp6454 = tmp4025 ? const_555_127 : tmp6373;
    assign tmp6506 = _ver_out_tmp_40 == tmp7898;
    assign tmp6514 = {tmp4703, tmp4703};
    assign tmp6515 = {tmp6514, tmp7882};
    assign tmp6516 = {tmp4110[8]};
    assign tmp6519 = tmp6515 + tmp4116;
    assign tmp6533 = tmp4128 ^ tmp5887;
    assign tmp6539 = {tmp4136[9]};
    assign tmp6542 = tmp6539 ^ tmp6140;
    assign tmp6544 = ~tmp6516;
    assign tmp6551 = tmp4119 - tmp5375;
    assign tmp6552 = {tmp6551[8]};
    assign tmp6555 = tmp6552 ^ tmp6597;
    assign tmp6566 = tmp7882 - tmp5375;
    assign tmp6567 = {tmp6566[8]};
    assign tmp6573 = tmp5888 ^ tmp1604;
    assign tmp6579 = {tmp4176[9]};
    assign tmp6597 = ~tmp4194;
    assign tmp6601 = tmp4184 & tmp4198;
    assign tmp6653 = ~tmp5986;
    assign tmp6665 = ~tmp2753;
    assign tmp6680 = tmp6356 & tmp6653;
    assign tmp6732 = tmp5375 - tmp10;
    assign tmp6738 = tmp7027 ? tmp7034 : tmp7036;
    assign tmp6740 = tmp1893 == const_581_1;
    assign tmp6753 = tmp6738 - tmp7053;
    assign tmp6754 = {tmp6753[9]};
    assign tmp6755 = {tmp6738[8]};
    assign tmp6756 = ~tmp6755;
    assign tmp6757 = tmp6754 ^ tmp6756;
    assign tmp6759 = ~tmp7061;
    assign tmp6760 = tmp6757 ^ tmp6759;
    assign tmp6761 = {tmp11[7]};
    assign tmp6762 = tmp6761 == const_588_1;
    assign tmp6763 = tmp11 == _ver_out_tmp_55;
    assign tmp6771 = {const_594_0, tmp11};
    assign tmp6772 = tmp6762 ? tmp2481 : tmp6771;
    assign tmp6774 = tmp349 == const_595_1;
    assign tmp6787 = tmp6772 - tmp7094;
    assign tmp6788 = {tmp6787[9]};
    assign tmp6789 = {tmp6772[8]};
    assign tmp6790 = ~tmp6789;
    assign tmp6791 = tmp6788 ^ tmp6790;
    assign tmp6792 = {tmp7094[8]};
    assign tmp6794 = tmp6791 ^ tmp7103;
    assign tmp6795 = tmp6760 & tmp6794;
    assign tmp6798 = tmp12 == _ver_out_tmp_61;
    assign tmp6816 = tmp7126 ? tmp4109 : tmp2573;
    assign tmp6818 = {const_615_0, tmp16};
    assign tmp6819 = tmp7125 ? tmp6816 : tmp6818;
    assign tmp6822 = tmp7119 - tmp6819;
    assign tmp6823 = {tmp6822[9]};
    assign tmp6824 = {tmp7119[8]};
    assign tmp6825 = ~tmp6824;
    assign tmp6826 = tmp6823 ^ tmp6825;
    assign tmp6828 = ~tmp7143;
    assign tmp6829 = tmp6826 ^ tmp6828;
    assign tmp6830 = tmp6795 & tmp6829;
    assign tmp6832 = tmp711 == const_616_1;
    assign tmp6841 = {const_622_0, tmp13};
    assign tmp6844 = tmp7579 == const_623_1;
    assign tmp6848 = tmp5375 - tmp17;
    assign tmp6853 = {const_629_0, tmp17};
    assign tmp6857 = tmp7160 - tmp7176;
    assign tmp6858 = {tmp6857[9]};
    assign tmp6859 = {tmp7160[8]};
    assign tmp6860 = ~tmp6859;
    assign tmp6861 = tmp6858 ^ tmp6860;
    assign tmp6862 = {tmp7176[8]};
    assign tmp6864 = tmp6861 ^ tmp7185;
    assign tmp6865 = tmp6830 & tmp6864;
    assign tmp6942 = ~tmp7865;
    assign tmp6951 = ~tmp79;
    assign tmp6991 = tmp7385 & tmp6942;
    assign tmp7009 = tmp6991 & tmp6865;
    assign tmp7026 = {tmp10[7]};
    assign tmp7027 = tmp7026 == const_632_1;
    assign tmp7034 = tmp2089 ? tmp4109 : tmp6732;
    assign tmp7036 = {const_638_0, tmp10};
    assign tmp7038 = {tmp6738[8], tmp6738[7], tmp6738[6], tmp6738[5], tmp6738[4], tmp6738[3], tmp6738[2], tmp6738[1]};
    assign tmp7039 = {tmp7038[7]};
    assign tmp7041 = {tmp7039, tmp7038};
    assign tmp7052 = {const_645_0, tmp14};
    assign tmp7053 = tmp6740 ? tmp1064 : tmp7052;
    assign tmp7056 = tmp7053 - tmp7041;
    assign tmp7057 = {tmp7056[9]};
    assign tmp7058 = {tmp7041[8]};
    assign tmp7059 = ~tmp7058;
    assign tmp7060 = tmp7057 ^ tmp7059;
    assign tmp7061 = {tmp7053[8]};
    assign tmp7063 = tmp7060 ^ tmp6759;
    assign tmp7064 = tmp7041 == tmp7053;
    assign tmp7065 = tmp7063 | tmp7064;
    assign tmp7066 = tmp18 & tmp7065;
    assign tmp7079 = {tmp6772[8], tmp6772[7], tmp6772[6], tmp6772[5], tmp6772[4], tmp6772[3], tmp6772[2], tmp6772[1]};
    assign tmp7080 = {tmp7079[7]};
    assign tmp7082 = {tmp7080, tmp7079};
    assign tmp7093 = {const_659_0, tmp15};
    assign tmp7094 = tmp6774 ? tmp1089 : tmp7093;
    assign tmp7097 = tmp7094 - tmp7082;
    assign tmp7098 = {tmp7097[9]};
    assign tmp7099 = {tmp7082[8]};
    assign tmp7100 = ~tmp7099;
    assign tmp7101 = tmp7098 ^ tmp7100;
    assign tmp7103 = ~tmp6792;
    assign tmp7104 = tmp7101 ^ tmp7103;
    assign tmp7105 = tmp7082 == tmp7094;
    assign tmp7106 = tmp7104 | tmp7105;
    assign tmp7107 = tmp7066 & tmp7106;
    assign tmp7109 = tmp1731 == const_660_1;
    assign tmp7118 = {const_666_0, tmp12};
    assign tmp7119 = tmp7109 ? tmp2500 : tmp7118;
    assign tmp7120 = {tmp7119[8], tmp7119[7], tmp7119[6], tmp7119[5], tmp7119[4], tmp7119[3], tmp7119[2], tmp7119[1]};
    assign tmp7121 = {tmp7120[7]};
    assign tmp7123 = {tmp7121, tmp7120};
    assign tmp7125 = tmp1396 == const_667_1;
    assign tmp7126 = tmp16 == _ver_out_tmp_2;
    assign tmp7138 = tmp6819 - tmp7123;
    assign tmp7139 = {tmp7138[9]};
    assign tmp7140 = {tmp7123[8]};
    assign tmp7141 = ~tmp7140;
    assign tmp7142 = tmp7139 ^ tmp7141;
    assign tmp7143 = {tmp6819[8]};
    assign tmp7145 = tmp7142 ^ tmp6828;
    assign tmp7146 = tmp7123 == tmp6819;
    assign tmp7147 = tmp7145 | tmp7146;
    assign tmp7148 = tmp7107 & tmp7147;
    assign tmp7151 = tmp13 == _ver_out_tmp_5;
    assign tmp7157 = tmp7151 ? tmp4109 : tmp2516;
    assign tmp7160 = tmp6832 ? tmp7157 : tmp6841;
    assign tmp7161 = {tmp7160[8], tmp7160[7], tmp7160[6], tmp7160[5], tmp7160[4], tmp7160[3], tmp7160[2], tmp7160[1]};
    assign tmp7162 = {tmp7161[7]};
    assign tmp7164 = {tmp7162, tmp7161};
    assign tmp7176 = tmp6844 ? tmp2595 : tmp6853;
    assign tmp7179 = tmp7176 - tmp7164;
    assign tmp7180 = {tmp7179[9]};
    assign tmp7181 = {tmp7164[8]};
    assign tmp7182 = ~tmp7181;
    assign tmp7183 = tmp7180 ^ tmp7182;
    assign tmp7185 = ~tmp6862;
    assign tmp7186 = tmp7183 ^ tmp7185;
    assign tmp7187 = tmp7164 == tmp7176;
    assign tmp7188 = tmp7186 | tmp7187;
    assign tmp7189 = tmp7148 & tmp7188;
    assign tmp7226 = {tmp10[7], tmp10[6], tmp10[5], tmp10[4], tmp10[3], tmp10[2], tmp10[1]};
    assign tmp7227 = {tmp7226[6]};
    assign tmp7229 = {tmp7227, tmp7226};
    assign tmp7249 = {tmp11[7], tmp11[6], tmp11[5], tmp11[4], tmp11[3], tmp11[2], tmp11[1]};
    assign tmp7250 = {tmp7249[6]};
    assign tmp7252 = {tmp7250, tmp7249};
    assign tmp7270 = tmp7390 & tmp7189;
    assign tmp7272 = {tmp12[7], tmp12[6], tmp12[5], tmp12[4], tmp12[3], tmp12[2], tmp12[1]};
    assign tmp7273 = {tmp7272[6]};
    assign tmp7275 = {tmp7273, tmp7272};
    assign tmp7291 = ~tmp6865;
    assign tmp7294 = tmp7270 & tmp7866;
    assign tmp7295 = {tmp13[7], tmp13[6], tmp13[5], tmp13[4], tmp13[3], tmp13[2], tmp13[1]};
    assign tmp7296 = {tmp7295[6]};
    assign tmp7298 = {tmp7296, tmp7295};
    assign tmp7319 = {tmp1316, const_690_0};
    assign tmp7324 = tmp5375 - tmp14;
    assign tmp7325 = {tmp7324[8]};
    assign tmp7336 = tmp7319 - tmp5375;
    assign tmp7340 = tmp1335 ^ tmp320;
    assign tmp7343 = tmp7340 ^ tmp1604;
    assign tmp7344 = tmp1858 & tmp7343;
    assign tmp7350 = {tmp2624[8]};
    assign tmp7353 = tmp7350 ^ tmp283;
    assign tmp7356 = tmp7353 ^ tmp1604;
    assign tmp7365 = tmp1360 ^ tmp1604;
    assign tmp7368 = tmp7365 ^ tmp320;
    assign tmp7369 = tmp5375 == tmp7319;
    assign tmp7370 = tmp7368 | tmp7369;
    assign tmp7371 = tmp7356 & tmp7370;
    assign tmp7385 = tmp2549 & tmp6665;
    assign tmp7390 = tmp6991 & tmp7291;
    assign tmp7393 = tmp7270 & tmp3387;
    assign tmp7394 = {tmp15[6], tmp15[5], tmp15[4], tmp15[3], tmp15[2], tmp15[1], tmp15[0]};
    assign tmp7401 = {tmp344[8]};
    assign tmp7413 = {tmp356[8]};
    assign tmp7416 = tmp7413 ^ tmp359;
    assign tmp7420 = tmp1870 & tmp363;
    assign tmp7425 = tmp15 - tmp5375;
    assign tmp7426 = {tmp7425[8]};
    assign tmp7437 = tmp5375 - tmp339;
    assign tmp7444 = tmp385 ^ tmp359;
    assign tmp7446 = tmp7444 | tmp389;
    assign tmp7449 = tmp391 ? _ver_out_tmp_11 : tmp392;
    assign tmp7470 = {tmp16[6], tmp16[5], tmp16[4], tmp16[3], tmp16[2], tmp16[1], tmp16[0]};
    assign tmp7483 = tmp1395 ^ tmp2019;
    assign tmp7488 = tmp1386 - tmp5375;
    assign tmp7489 = {tmp7488[8]};
    assign tmp7492 = tmp7489 ^ tmp1434;
    assign tmp7495 = tmp7492 ^ tmp1604;
    assign tmp7496 = tmp7483 & tmp7495;
    assign tmp7508 = tmp1420 ^ tmp1604;
    assign tmp7520 = tmp1432 ^ tmp1434;
    assign tmp7523 = tmp7508 & tmp1437;
    assign tmp7525 = tmp7523 ? _ver_out_tmp_12 : tmp1439;
    assign tmp7546 = {tmp17[6], tmp17[5], tmp17[4], tmp17[3], tmp17[2], tmp17[1], tmp17[0]};
    assign tmp7547 = {tmp7546, const_711_0};
    assign tmp7553 = {tmp6848[8]};
    assign tmp7556 = tmp7553 ^ tmp1604;
    assign tmp7558 = ~tmp7579;
    assign tmp7564 = tmp7547 - tmp5375;
    assign tmp7565 = {tmp7564[8]};
    assign tmp7567 = ~tmp7594;
    assign tmp7568 = tmp7565 ^ tmp7567;
    assign tmp7571 = tmp7568 ^ tmp1604;
    assign tmp7572 = tmp918 & tmp7571;
    assign tmp7579 = {tmp17[7]};
    assign tmp7581 = tmp2355 ^ tmp7558;
    assign tmp7584 = tmp7581 ^ tmp1604;
    assign tmp7589 = tmp5375 - tmp7547;
    assign tmp7590 = {tmp7589[8]};
    assign tmp7593 = tmp7590 ^ tmp1604;
    assign tmp7594 = {tmp7547[7]};
    assign tmp7596 = tmp7593 ^ tmp7567;
    assign tmp7597 = tmp5375 == tmp7547;
    assign tmp7598 = tmp7596 | tmp7597;
    assign tmp7599 = tmp7584 & tmp7598;
    assign tmp7600 = tmp7572 ? const_716_127 : tmp7547;
    assign tmp7601 = tmp7599 ? _ver_out_tmp_13 : tmp7600;
    assign tmp7639 = ~tmp7189;
    assign tmp7640 = tmp7390 & tmp7639;
    assign tmp7692 = tmp68 ? const_6_0 : tmp10;
    assign tmp7693 = tmp337 ? tmp192 : tmp7692;
    assign tmp7694 = tmp489 ? tmp12 : tmp7693;
    assign tmp7695 = tmp1006 ? tmp613 : tmp7694;
    assign tmp7696 = tmp1107 ? tmp1015 : tmp7695;
    assign tmp7697 = tmp1384 ? tmp192 : tmp7696;
    assign tmp7698 = tmp1580 ? tmp11 : tmp7697;
    assign tmp7699 = tmp1820 ? tmp1678 : tmp7698;
    assign tmp7700 = tmp2169 ? tmp1015 : tmp7699;
    assign tmp7701 = tmp2895 ? tmp1015 : tmp7700;
    assign tmp7702 = tmp3079 ? tmp2921 : tmp7701;
    assign tmp7703 = tmp3222 ? tmp7870 : tmp7702;
    assign tmp7704 = tmp3701 ? tmp7886 : tmp7703;
    assign tmp7705 = tmp4362 ? tmp7886 : tmp7704;
    assign tmp7706 = tmp4931 ? tmp2921 : tmp7705;
    assign tmp7707 = tmp5077 ? tmp7870 : tmp7706;
    assign tmp7708 = tmp6209 ? tmp7886 : tmp7707;
    assign tmp7709 = tmp7009 ? tmp14 : tmp7708;
    assign tmp7710 = tmp7294 ? tmp7229 : tmp7709;
    assign tmp7711 = tmp68 ? const_7_2 : tmp11;
    assign tmp7712 = tmp337 ? tmp259 : tmp7711;
    assign tmp7713 = tmp489 ? tmp13 : tmp7712;
    assign tmp7714 = tmp1006 ? tmp734 : tmp7713;
    assign tmp7715 = tmp1107 ? tmp2482 : tmp7714;
    assign tmp7716 = tmp1133 ? tmp10 : tmp7715;
    assign tmp7717 = tmp1580 ? tmp10 : tmp7716;
    assign tmp7718 = tmp1820 ? tmp10 : tmp7717;
    assign tmp7719 = tmp2895 ? tmp2482 : tmp7718;
    assign tmp7720 = tmp3079 ? tmp2937 : tmp7719;
    assign tmp7721 = tmp3222 ? tmp7874 : tmp7720;
    assign tmp7722 = tmp3701 ? tmp7890 : tmp7721;
    assign tmp7723 = tmp4362 ? tmp7890 : tmp7722;
    assign tmp7724 = tmp4931 ? tmp2937 : tmp7723;
    assign tmp7725 = tmp5077 ? tmp7874 : tmp7724;
    assign tmp7726 = tmp6209 ? tmp7890 : tmp7725;
    assign tmp7727 = tmp7009 ? tmp15 : tmp7726;
    assign tmp7728 = tmp7294 ? tmp7252 : tmp7727;
    assign tmp7729 = tmp68 ? const_8_1 : tmp12;
    assign tmp7730 = tmp107 ? tmp10 : tmp7729;
    assign tmp7731 = tmp489 ? tmp10 : tmp7730;
    assign tmp7732 = tmp1006 ? tmp10 : tmp7731;
    assign tmp7733 = tmp1384 ? tmp1302 : tmp7732;
    assign tmp7734 = tmp1580 ? tmp13 : tmp7733;
    assign tmp7735 = tmp1820 ? tmp1803 : tmp7734;
    assign tmp7736 = tmp2169 ? tmp2501 : tmp7735;
    assign tmp7737 = tmp2895 ? tmp2501 : tmp7736;
    assign tmp7738 = tmp3079 ? tmp3062 : tmp7737;
    assign tmp7739 = tmp3222 ? tmp7878 : tmp7738;
    assign tmp7740 = tmp3701 ? tmp7894 : tmp7739;
    assign tmp7741 = tmp4362 ? tmp7894 : tmp7740;
    assign tmp7742 = tmp4931 ? tmp3062 : tmp7741;
    assign tmp7743 = tmp5077 ? tmp7878 : tmp7742;
    assign tmp7744 = tmp6209 ? tmp7894 : tmp7743;
    assign tmp7745 = tmp7009 ? tmp16 : tmp7744;
    assign tmp7746 = tmp7294 ? tmp7275 : tmp7745;
    assign tmp7747 = tmp68 ? const_9_0 : tmp13;
    assign tmp7748 = tmp107 ? tmp11 : tmp7747;
    assign tmp7749 = tmp489 ? tmp11 : tmp7748;
    assign tmp7750 = tmp1006 ? tmp11 : tmp7749;
    assign tmp7751 = tmp1133 ? tmp12 : tmp7750;
    assign tmp7752 = tmp1580 ? tmp12 : tmp7751;
    assign tmp7753 = tmp1820 ? tmp12 : tmp7752;
    assign tmp7754 = tmp2895 ? tmp2520 : tmp7753;
    assign tmp7755 = tmp3079 ? tmp3083 : tmp7754;
    assign tmp7756 = tmp3222 ? tmp7882 : tmp7755;
    assign tmp7757 = tmp3701 ? tmp7898 : tmp7756;
    assign tmp7758 = tmp4362 ? tmp7898 : tmp7757;
    assign tmp7759 = tmp4931 ? tmp3083 : tmp7758;
    assign tmp7760 = tmp5077 ? tmp7882 : tmp7759;
    assign tmp7761 = tmp6209 ? tmp7898 : tmp7760;
    assign tmp7762 = tmp7009 ? tmp17 : tmp7761;
    assign tmp7763 = tmp7294 ? tmp7298 : tmp7762;
    assign tmp7764 = tmp68 ? const_10_0 : tmp14;
    assign tmp7765 = tmp337 ? tmp326 : tmp7764;
    assign tmp7766 = tmp489 ? tmp16 : tmp7765;
    assign tmp7767 = tmp1006 ? tmp855 : tmp7766;
    assign tmp7768 = tmp1107 ? tmp2539 : tmp7767;
    assign tmp7769 = tmp1384 ? tmp326 : tmp7768;
    assign tmp7770 = tmp1580 ? tmp15 : tmp7769;
    assign tmp7771 = tmp1820 ? tmp1928 : tmp7770;
    assign tmp7772 = tmp2169 ? tmp2539 : tmp7771;
    assign tmp7773 = tmp3079 ? tmp7886 : tmp7772;
    assign tmp7774 = tmp3222 ? tmp5183 : tmp7773;
    assign tmp7775 = tmp3701 ? tmp3799 : tmp7774;
    assign tmp7776 = tmp4362 ? tmp7870 : tmp7775;
    assign tmp7777 = tmp4931 ? tmp7886 : tmp7776;
    assign tmp7778 = tmp5077 ? tmp5183 : tmp7777;
    assign tmp7779 = tmp6209 ? tmp3799 : tmp7778;
    assign tmp7780 = tmp7009 ? tmp10 : tmp7779;
    assign tmp7781 = tmp7393 ? tmp326 : tmp7780;
    assign tmp7782 = tmp68 ? const_11_0 : tmp15;
    assign tmp7783 = tmp337 ? tmp7449 : tmp7782;
    assign tmp7784 = tmp489 ? tmp17 : tmp7783;
    assign tmp7785 = tmp1006 ? tmp976 : tmp7784;
    assign tmp7786 = tmp1107 ? tmp2558 : tmp7785;
    assign tmp7787 = tmp1133 ? tmp14 : tmp7786;
    assign tmp7788 = tmp1580 ? tmp14 : tmp7787;
    assign tmp7789 = tmp1820 ? tmp14 : tmp7788;
    assign tmp7790 = tmp3079 ? tmp7890 : tmp7789;
    assign tmp7791 = tmp3222 ? tmp3370 : tmp7790;
    assign tmp7792 = tmp3701 ? tmp3933 : tmp7791;
    assign tmp7793 = tmp4362 ? tmp7874 : tmp7792;
    assign tmp7794 = tmp4931 ? tmp7890 : tmp7793;
    assign tmp7795 = tmp5077 ? tmp3370 : tmp7794;
    assign tmp7796 = tmp6209 ? tmp3933 : tmp7795;
    assign tmp7797 = tmp7009 ? tmp11 : tmp7796;
    assign tmp7798 = tmp7393 ? tmp7449 : tmp7797;
    assign tmp7799 = tmp68 ? const_12_0 : tmp16;
    assign tmp7800 = tmp107 ? tmp14 : tmp7799;
    assign tmp7801 = tmp489 ? tmp14 : tmp7800;
    assign tmp7802 = tmp1006 ? tmp14 : tmp7801;
    assign tmp7803 = tmp1384 ? tmp7525 : tmp7802;
    assign tmp7804 = tmp1580 ? tmp17 : tmp7803;
    assign tmp7805 = tmp1820 ? tmp2053 : tmp7804;
    assign tmp7806 = tmp2169 ? tmp2577 : tmp7805;
    assign tmp7807 = tmp3079 ? tmp7894 : tmp7806;
    assign tmp7808 = tmp3222 ? tmp3444 : tmp7807;
    assign tmp7809 = tmp3701 ? tmp4067 : tmp7808;
    assign tmp7810 = tmp4362 ? tmp7878 : tmp7809;
    assign tmp7811 = tmp4931 ? tmp7894 : tmp7810;
    assign tmp7812 = tmp5077 ? tmp3444 : tmp7811;
    assign tmp7813 = tmp6209 ? tmp4067 : tmp7812;
    assign tmp7814 = tmp7009 ? tmp12 : tmp7813;
    assign tmp7815 = tmp7393 ? tmp7525 : tmp7814;
    assign tmp7816 = tmp68 ? const_13_1 : tmp17;
    assign tmp7817 = tmp107 ? tmp15 : tmp7816;
    assign tmp7818 = tmp489 ? tmp15 : tmp7817;
    assign tmp7819 = tmp1006 ? tmp15 : tmp7818;
    assign tmp7820 = tmp1133 ? tmp16 : tmp7819;
    assign tmp7821 = tmp1580 ? tmp16 : tmp7820;
    assign tmp7822 = tmp1820 ? tmp16 : tmp7821;
    assign tmp7823 = tmp3079 ? tmp7898 : tmp7822;
    assign tmp7824 = tmp3222 ? tmp3518 : tmp7823;
    assign tmp7825 = tmp3701 ? tmp4201 : tmp7824;
    assign tmp7826 = tmp4362 ? tmp7882 : tmp7825;
    assign tmp7827 = tmp4931 ? tmp7898 : tmp7826;
    assign tmp7828 = tmp5077 ? tmp3518 : tmp7827;
    assign tmp7829 = tmp6209 ? tmp4201 : tmp7828;
    assign tmp7830 = tmp7009 ? tmp13 : tmp7829;
    assign tmp7831 = tmp7393 ? tmp7601 : tmp7830;
    assign tmp7832 = tmp68 ? const_14_0 : tmp18;
    assign tmp7833 = tmp997 ? tmp18 : tmp7832;
    assign tmp7834 = tmp1953 ? tmp18 : tmp7833;
    assign tmp7835 = tmp2764 ? const_291_0 : tmp7834;
    assign tmp7836 = tmp2895 ? const_295_0 : tmp7835;
    assign tmp7837 = tmp3150 ? const_317_0 : tmp7836;
    assign tmp7838 = tmp3701 ? const_347_0 : tmp7837;
    assign tmp7839 = tmp4362 ? const_401_0 : tmp7838;
    assign tmp7840 = tmp4796 ? const_431_0 : tmp7839;
    assign tmp7841 = tmp6209 ? const_517_1 : tmp7840;
    assign tmp7842 = tmp6680 ? const_571_0 : tmp7841;
    assign tmp7843 = const_758_0 ? const_573_0 : tmp7842;
    assign tmp7844 = tmp7009 ? const_631_1 : tmp7843;
    assign tmp7845 = tmp7270 ? const_689_1 : tmp7844;
    assign tmp7846 = tmp7640 ? tmp18 : tmp7845;
    assign tmp7847 = const_759_0 ? tmp18 : tmp7846;
    assign tmp7848 = tmp68 ? const_15_0 : my_calculator_out_z;
    assign tmp7849 = tmp2764 ? const_290_15 : tmp7848;
    assign tmp7850 = tmp2895 ? const_294_8 : tmp7849;
    assign tmp7851 = tmp3150 ? const_316_1 : tmp7850;
    assign tmp7852 = tmp3701 ? const_346_4 : tmp7851;
    assign tmp7853 = tmp4362 ? const_400_6 : tmp7852;
    assign tmp7854 = tmp4796 ? const_430_2 : tmp7853;
    assign tmp7855 = tmp6209 ? const_516_5 : tmp7854;
    assign tmp7856 = tmp6680 ? const_570_0 : tmp7855;
    assign tmp7857 = const_757_0 ? const_572_0 : tmp7856;
    assign tmp7858 = tmp7009 ? const_630_7 : tmp7857;
    assign tmp7859 = tmp7270 ? const_688_3 : tmp7858;
    assign tmp7860 = tmp7640 ? const_718_0 : tmp7859;
    assign tmp7861 = const_756_0 ? const_719_0 : tmp7860;
    assign tmp7862 = tmp2549 ? tmp2276 : const_720_0;
    assign tmp7863 = tmp2549 ? tmp2363 : const_721_0;
    assign tmp7864 = tmp2549 ? tmp2388 : const_722_0;
    assign tmp7865 = tmp2549 ? tmp2401 : const_723_0;
    assign tmp7866 = tmp2549 ? tmp2419 : const_724_0;
    assign tmp7869 = tmp2512 ? tmp1015 : tmp5375;
    assign tmp7870 = tmp2660 ? tmp10 : tmp7869;
    assign tmp7873 = tmp2512 ? tmp2482 : tmp5375;
    assign tmp7874 = tmp2660 ? tmp11 : tmp7873;
    assign tmp7877 = tmp2512 ? tmp2501 : tmp5375;
    assign tmp7878 = tmp2660 ? tmp12 : tmp7877;
    assign tmp7881 = tmp2512 ? tmp2520 : tmp5375;
    assign tmp7882 = tmp2660 ? tmp13 : tmp7881;
    assign tmp7885 = tmp2512 ? tmp2539 : tmp5375;
    assign tmp7886 = tmp2660 ? tmp14 : tmp7885;
    assign tmp7889 = tmp2512 ? tmp2558 : tmp5375;
    assign tmp7890 = tmp2660 ? tmp15 : tmp7889;
    assign tmp7893 = tmp2512 ? tmp2577 : tmp5375;
    assign tmp7894 = tmp2660 ? tmp16 : tmp7893;
    assign tmp7897 = tmp2512 ? tmp2596 : tmp5375;
    assign tmp7898 = tmp2660 ? tmp17 : tmp7897;
    assign tmp7908 = my_calculator_out_z == tmp87;
    assign tmp7914 = my_calculator_out_z == tmp127;
    assign tmp7917 = my_calculator_out_z == tmp517;
    assign tmp7918 = tmp7914 | tmp7917;
    assign tmp7919 = my_calculator_out_z == const_749_15;
    assign tmp7920 = tmp7918 | tmp7919;
    assign tmp7921 = {tmp0[25]};
    assign tmp7923 = ~tmp8;
    assign tmp7924 = {const_751_0, const_751_0, const_751_0, const_751_0};
    assign tmp7925 = {tmp7924, const_750_1};
    assign tmp7926 = tmp7899 + tmp7925;
    assign tmp7927 = {tmp7926[4], tmp7926[3], tmp7926[2], tmp7926[1], tmp7926[0]};
    assign tmp7928 = tmp7923 ? tmp7927 : tmp7899;

    // Registers
    always @(posedge clk)
    begin
        begin
            my_calculator_ctrl <= tmp7903;
            my_calculator_in_x <= tmp7904;
            my_calculator_in_y <= tmp7905;
            my_calculator_out_z <= tmp7861;
            tmp0 <= tmp4;
            tmp5 <= tmp7921;
            tmp10 <= tmp7710;
            tmp11 <= tmp7728;
            tmp12 <= tmp7746;
            tmp13 <= tmp7763;
            tmp14 <= tmp7781;
            tmp15 <= tmp7798;
            tmp16 <= tmp7815;
            tmp17 <= tmp7831;
            tmp18 <= tmp7847;
            tmp7899 <= tmp7928;
            was_toggled <= tmp7923;
        end
    end

    // Memory mem_0: tmp7900
    assign tmp7903 = mem_0[tmp7899];

    // Memory mem_1: tmp7901
    assign tmp7904 = mem_1[tmp7899];

    // Memory mem_2: tmp7902
    assign tmp7905 = mem_2[tmp7899];

endmodule

