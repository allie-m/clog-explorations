// Simple tri-colour LED blink example.

// Correctly map pins for the iCE40UP5K SB_RGBA_DRV hard macro.

`define GREENPWM RGB0PWM
`define REDPWM   RGB1PWM
`define BLUEPWM  RGB2PWM

// taken (mostly) from
// https://github.com/im-tomu/fomu-workshop/blob/master/hdl/verilog/blink-expanded/blink.v

module top (
    // 48MHz Clock input
    // --------
    input clki,
    // LED outputs
    // --------
    output rgb0,
    output rgb1,
    output rgb2,
    // User touchable pins
    // --------
    // Connect 1-2 to enable blue LED
    input  user_1,
    output user_2,
    // Connect 3-4 to enable red LED
    output user_3,
    input  user_4,
    // USB Pins (which should be statically driven if not being used).
    // --------
    output usb_dp,
    output usb_dn,
    output usb_dp_pu
);

    // Assign USB pins to "0" so as to disconnect Fomu from
    // the host system.  Otherwise it would try to talk to
    // us over USB, which wouldn't work since we have no stack.
    assign usb_dp = 1'b0;
    assign usb_dn = 1'b0;
    assign usb_dp_pu = 1'b0;
    // Configure user pins so that we can detect the user connecting
    // 1-2 or 3-4 with conductive material.
    //
    // We do this by grounding user_2 and user_3, and configuring inputs
    // with pullups on user_1 and user_4.
    assign user_2 = 1'b0;
    assign user_3 = 1'b0;

    // Connect to system clock (with buffering)
    wire clk;
    SB_GB clk_gb (
        .USER_SIGNAL_TO_GLOBAL_BUFFER(clki),
        .GLOBAL_BUFFER_OUTPUT(clk)
    );

    // PyRTL module goes here:
    wire [3:0] colors;
    toplevel pyrtl_toplevel (
        .clk (clk),
        .in_1 (~user_1),
        .in_2 (~user_4),
        .red_o (colors[0]),
        .green_o (colors[1]),
        .blue_o (colors[2])
    );

    // Instantiate iCE40 LED driver hard logic, connecting up
    // counter state and LEDs.
    //
    // Note that it's possible to drive the LEDs directly,
    // however that is not current-limited and results in
    // overvolting the red LED.
    //
    // See also:
    // https://www.latticesemi.com/-/media/LatticeSemi/Documents/ApplicationNotes/IK/ICE40LEDDriverUsageGuide.ashx?document_id=50668
    SB_RGBA_DRV #(
        .CURRENT_MODE("0b1"),       // half current
        .RGB0_CURRENT("0b000011"),  // 4 mA
        .RGB1_CURRENT("0b000011"),  // 4 mA
        .RGB2_CURRENT("0b000011")   // 4 mA
    ) RGBA_DRIVER (
        .CURREN(1'b1),
        .RGBLEDEN(1'b1),
        .`REDPWM(colors[0]),      // Red
        .`GREENPWM(colors[1]),    // Green
        .`BLUEPWM(colors[2]),     // Blue
        .RGB0(rgb0),
        .RGB1(rgb1),
        .RGB2(rgb2)
    );

endmodule
// Generated automatically via PyRTL
// As one initial test of synthesis, map to FPGA with:
//   yosys -p "synth_xilinx -top toplevel" thisfile.v

module toplevel(clk, in_1, in_2, blue_o, green_o, red_o);
    input clk;
    input in_1;
    input in_2;
    output blue_o;
    output green_o;
    output red_o;

    reg[25:0] tmp0;
    reg tmp5;
    reg tmp7;
    reg[255:0] tmp11;
    reg[255:0] tmp12;
    reg[255:0] tmp13;
    reg[255:0] tmp14;
    reg[255:0] tmp15;
    reg[255:0] tmp16;
    reg[255:0] tmp17;
    reg[255:0] tmp18;
    reg tmp19;
    reg[2:0] tmp7688;

    wire[255:0] _ver_out_tmp_0;
    wire[255:0] _ver_out_tmp_1;
    wire[255:0] _ver_out_tmp_2;
    wire[255:0] _ver_out_tmp_3;
    wire[255:0] _ver_out_tmp_4;
    wire[255:0] _ver_out_tmp_5;
    wire[255:0] _ver_out_tmp_6;
    wire[255:0] _ver_out_tmp_7;
    wire[255:0] _ver_out_tmp_8;
    wire[255:0] _ver_out_tmp_9;
    wire[255:0] _ver_out_tmp_10;
    wire[255:0] _ver_out_tmp_11;
    wire[255:0] _ver_out_tmp_12;
    wire[255:0] _ver_out_tmp_13;
    wire[255:0] _ver_out_tmp_14;
    wire[255:0] _ver_out_tmp_15;
    wire[255:0] _ver_out_tmp_16;
    wire[255:0] _ver_out_tmp_17;
    wire[255:0] _ver_out_tmp_18;
    wire[255:0] _ver_out_tmp_19;
    wire[255:0] _ver_out_tmp_20;
    wire[255:0] _ver_out_tmp_21;
    wire[255:0] _ver_out_tmp_22;
    wire[255:0] _ver_out_tmp_23;
    wire[255:0] _ver_out_tmp_24;
    wire[255:0] _ver_out_tmp_25;
    wire[255:0] _ver_out_tmp_26;
    wire[255:0] _ver_out_tmp_27;
    wire[255:0] _ver_out_tmp_28;
    wire[255:0] _ver_out_tmp_29;
    wire[255:0] _ver_out_tmp_30;
    wire[255:0] _ver_out_tmp_31;
    wire[255:0] _ver_out_tmp_32;
    wire[255:0] _ver_out_tmp_33;
    wire[255:0] _ver_out_tmp_34;
    wire[255:0] _ver_out_tmp_35;
    wire[255:0] _ver_out_tmp_36;
    wire[255:0] _ver_out_tmp_37;
    wire[255:0] _ver_out_tmp_38;
    wire[255:0] _ver_out_tmp_39;
    wire[255:0] _ver_out_tmp_40;
    wire[255:0] _ver_out_tmp_41;
    wire[255:0] _ver_out_tmp_42;
    wire[255:0] _ver_out_tmp_43;
    wire[255:0] _ver_out_tmp_44;
    wire[255:0] _ver_out_tmp_45;
    wire[255:0] _ver_out_tmp_46;
    wire[255:0] _ver_out_tmp_47;
    wire[255:0] _ver_out_tmp_48;
    wire[255:0] _ver_out_tmp_49;
    wire[255:0] _ver_out_tmp_50;
    wire[255:0] _ver_out_tmp_51;
    wire[255:0] _ver_out_tmp_52;
    wire[255:0] _ver_out_tmp_53;
    wire[255:0] _ver_out_tmp_54;
    wire[255:0] _ver_out_tmp_55;
    wire[255:0] _ver_out_tmp_56;
    wire[255:0] _ver_out_tmp_57;
    wire[255:0] _ver_out_tmp_58;
    wire[255:0] _ver_out_tmp_59;
    wire[255:0] _ver_out_tmp_60;
    wire[255:0] _ver_out_tmp_61;
    wire[255:0] _ver_out_tmp_62;
    wire[255:0] _ver_out_tmp_63;
    wire[255:0] _ver_out_tmp_64;
    wire[255:0] _ver_out_tmp_65;
    wire[255:0] _ver_out_tmp_66;
    wire[255:0] _ver_out_tmp_67;
    wire[255:0] _ver_out_tmp_68;
    wire[255:0] _ver_out_tmp_69;
    wire[255:0] _ver_out_tmp_70;
    wire[255:0] _ver_out_tmp_71;
    wire[255:0] _ver_out_tmp_72;
    wire[255:0] _ver_out_tmp_73;
    wire[255:0] _ver_out_tmp_74;
    wire[255:0] _ver_out_tmp_75;
    wire[255:0] _ver_out_tmp_76;
    wire[255:0] _ver_out_tmp_77;
    wire[255:0] _ver_out_tmp_78;
    wire[255:0] _ver_out_tmp_79;
    wire[255:0] _ver_out_tmp_80;
    wire[255:0] _ver_out_tmp_81;
    wire[255:0] _ver_out_tmp_82;
    wire[255:0] _ver_out_tmp_83;
    wire[255:0] _ver_out_tmp_84;
    wire[255:0] _ver_out_tmp_85;
    wire[255:0] _ver_out_tmp_86;
    wire[255:0] _ver_out_tmp_87;
    wire[255:0] _ver_out_tmp_88;
    wire[255:0] _ver_out_tmp_89;
    wire[255:0] _ver_out_tmp_90;
    wire[255:0] _ver_out_tmp_91;
    wire cfg_speculative_egest;
    wire const_0_1;
    wire const_1_1;
    wire const_2_0;
    wire const_3_0;
    wire const_4_0;
    wire[2:0] const_5_4;
    wire[255:0] const_6_0;
    wire[255:0] const_7_2;
    wire[255:0] const_8_1;
    wire[255:0] const_9_0;
    wire[255:0] const_10_0;
    wire[255:0] const_11_0;
    wire[255:0] const_12_0;
    wire[255:0] const_13_1;
    wire const_14_0;
    wire const_15_1;
    wire const_16_0;
    wire[3:0] const_17_0;
    wire const_18_0;
    wire const_19_0;
    wire[3:0] const_20_15;
    wire const_21_1;
    wire const_22_0;
    wire[1:0] const_23_2;
    wire const_24_0;
    wire[1:0] const_25_3;
    wire const_26_0;
    wire const_27_0;
    wire const_28_0;
    wire const_29_0;
    wire const_30_0;
    wire const_31_0;
    wire[255:0] const_32_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_34_0;
    wire const_35_0;
    wire const_36_0;
    wire const_37_0;
    wire const_38_0;
    wire[255:0] const_39_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_41_0;
    wire const_42_0;
    wire const_43_0;
    wire const_44_0;
    wire const_45_0;
    wire[255:0] const_46_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_48_0;
    wire const_49_0;
    wire const_50_0;
    wire const_51_0;
    wire const_52_0;
    wire[255:0] const_53_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire[2:0] const_55_6;
    wire const_56_0;
    wire[2:0] const_57_7;
    wire const_58_0;
    wire[2:0] const_59_4;
    wire const_60_0;
    wire[2:0] const_61_5;
    wire const_62_0;
    wire const_63_0;
    wire const_64_0;
    wire const_65_0;
    wire const_66_0;
    wire const_67_0;
    wire const_68_0;
    wire[255:0] const_69_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_71_0;
    wire const_72_0;
    wire const_73_0;
    wire const_74_0;
    wire const_75_0;
    wire const_76_0;
    wire[255:0] const_77_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_79_0;
    wire const_80_0;
    wire const_81_0;
    wire const_82_0;
    wire const_83_0;
    wire const_84_0;
    wire[255:0] const_85_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_87_0;
    wire const_88_0;
    wire const_89_0;
    wire const_90_0;
    wire const_91_0;
    wire const_92_0;
    wire[255:0] const_93_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire[3:0] const_95_8;
    wire const_97_0;
    wire const_98_0;
    wire[254:0] const_99_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_100_0;
    wire const_102_0;
    wire const_103_0;
    wire[254:0] const_104_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_105_0;
    wire const_107_0;
    wire const_108_0;
    wire[254:0] const_109_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_110_0;
    wire const_112_0;
    wire const_113_0;
    wire[254:0] const_114_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_115_0;
    wire[1:0] const_116_2;
    wire const_117_0;
    wire[3:0] const_118_0;
    wire const_119_0;
    wire const_120_0;
    wire[3:0] const_121_15;
    wire const_122_1;
    wire const_123_0;
    wire[1:0] const_124_2;
    wire const_125_0;
    wire[1:0] const_126_3;
    wire const_127_0;
    wire const_128_0;
    wire const_129_0;
    wire const_130_0;
    wire const_131_0;
    wire const_132_0;
    wire[255:0] const_133_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_135_0;
    wire const_136_0;
    wire const_137_0;
    wire const_138_0;
    wire const_139_0;
    wire[255:0] const_140_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_142_0;
    wire const_143_0;
    wire const_144_0;
    wire const_145_0;
    wire const_146_0;
    wire[255:0] const_147_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_149_0;
    wire const_150_0;
    wire const_151_0;
    wire const_152_0;
    wire const_153_0;
    wire[255:0] const_154_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire[2:0] const_156_6;
    wire const_157_0;
    wire[2:0] const_158_7;
    wire const_159_0;
    wire[2:0] const_160_4;
    wire const_161_0;
    wire[2:0] const_162_5;
    wire const_163_0;
    wire const_164_0;
    wire const_165_0;
    wire const_166_0;
    wire const_167_0;
    wire const_168_0;
    wire const_169_0;
    wire[255:0] const_170_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_172_0;
    wire const_173_0;
    wire const_174_0;
    wire const_175_0;
    wire const_176_0;
    wire const_177_0;
    wire[255:0] const_178_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_180_0;
    wire const_181_0;
    wire const_182_0;
    wire const_183_0;
    wire const_184_0;
    wire const_185_0;
    wire[255:0] const_186_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_188_0;
    wire const_189_0;
    wire const_190_0;
    wire const_191_0;
    wire const_192_0;
    wire const_193_0;
    wire[255:0] const_194_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire[3:0] const_196_8;
    wire const_198_0;
    wire const_199_0;
    wire[254:0] const_200_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_201_0;
    wire const_203_0;
    wire const_204_0;
    wire[254:0] const_205_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_206_0;
    wire const_208_0;
    wire const_209_0;
    wire[254:0] const_210_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_211_0;
    wire const_213_0;
    wire const_214_0;
    wire[254:0] const_215_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_216_0;
    wire[1:0] const_217_3;
    wire const_218_0;
    wire const_219_0;
    wire const_220_0;
    wire const_221_0;
    wire const_222_0;
    wire const_223_0;
    wire const_224_0;
    wire const_225_0;
    wire const_226_0;
    wire const_227_0;
    wire const_228_0;
    wire const_229_0;
    wire const_230_0;
    wire const_231_0;
    wire const_232_0;
    wire const_233_0;
    wire const_234_0;
    wire const_235_0;
    wire const_236_0;
    wire const_237_0;
    wire const_238_0;
    wire const_239_0;
    wire const_240_0;
    wire const_242_0;
    wire const_243_0;
    wire[254:0] const_244_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_245_0;
    wire const_247_0;
    wire const_248_0;
    wire[254:0] const_249_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_250_0;
    wire const_252_0;
    wire const_253_0;
    wire[254:0] const_254_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_255_0;
    wire const_257_0;
    wire const_258_0;
    wire[254:0] const_259_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_260_0;
    wire const_262_0;
    wire const_263_0;
    wire[254:0] const_264_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_265_0;
    wire const_267_0;
    wire const_268_0;
    wire[254:0] const_269_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_270_0;
    wire const_272_0;
    wire const_273_0;
    wire[254:0] const_274_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_275_0;
    wire const_277_0;
    wire const_278_0;
    wire[254:0] const_279_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_280_0;
    wire const_281_0;
    wire const_282_0;
    wire const_283_0;
    wire const_284_0;
    wire const_285_0;
    wire const_286_0;
    wire const_287_0;
    wire const_288_0;
    wire const_289_0;
    wire const_290_0;
    wire[3:0] const_291_15;
    wire const_292_0;
    wire const_293_0;
    wire const_294_0;
    wire[3:0] const_295_8;
    wire const_296_0;
    wire const_298_0;
    wire const_299_0;
    wire[254:0] const_300_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_301_0;
    wire const_303_0;
    wire const_304_0;
    wire[254:0] const_305_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_306_0;
    wire const_308_0;
    wire const_309_0;
    wire[254:0] const_310_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_311_0;
    wire const_313_0;
    wire const_314_0;
    wire[254:0] const_315_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_316_0;
    wire[3:0] const_317_1;
    wire const_318_0;
    wire const_319_0;
    wire const_320_0;
    wire const_321_0;
    wire const_322_0;
    wire const_323_0;
    wire[255:0] const_324_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_326_0;
    wire const_327_0;
    wire const_328_0;
    wire const_329_0;
    wire const_330_0;
    wire[255:0] const_331_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_333_0;
    wire const_334_0;
    wire const_335_0;
    wire const_336_0;
    wire const_337_0;
    wire[255:0] const_338_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_340_0;
    wire const_341_0;
    wire const_342_0;
    wire const_343_0;
    wire const_344_0;
    wire[255:0] const_345_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire[3:0] const_347_4;
    wire const_348_0;
    wire const_350_0;
    wire const_351_0;
    wire[254:0] const_352_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_353_0;
    wire const_354_0;
    wire const_355_0;
    wire const_356_0;
    wire const_357_0;
    wire const_358_0;
    wire const_359_0;
    wire[255:0] const_360_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_363_0;
    wire const_364_0;
    wire[254:0] const_365_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_366_0;
    wire const_367_0;
    wire const_368_0;
    wire const_369_0;
    wire const_370_0;
    wire const_371_0;
    wire const_372_0;
    wire[255:0] const_373_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_376_0;
    wire const_377_0;
    wire[254:0] const_378_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_379_0;
    wire const_380_0;
    wire const_381_0;
    wire const_382_0;
    wire const_383_0;
    wire const_384_0;
    wire const_385_0;
    wire[255:0] const_386_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_389_0;
    wire const_390_0;
    wire[254:0] const_391_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_392_0;
    wire const_393_0;
    wire const_394_0;
    wire const_395_0;
    wire const_396_0;
    wire const_397_0;
    wire const_398_0;
    wire[255:0] const_399_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire[3:0] const_401_6;
    wire const_402_0;
    wire[1:0] const_403_0;
    wire const_404_0;
    wire const_405_0;
    wire const_406_0;
    wire const_407_0;
    wire[255:0] const_408_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire[1:0] const_410_0;
    wire const_411_0;
    wire const_412_0;
    wire const_413_0;
    wire const_414_0;
    wire[255:0] const_415_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire[1:0] const_417_0;
    wire const_418_0;
    wire const_419_0;
    wire const_420_0;
    wire const_421_0;
    wire[255:0] const_422_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire[1:0] const_424_0;
    wire const_425_0;
    wire const_426_0;
    wire const_427_0;
    wire const_428_0;
    wire[255:0] const_429_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire[3:0] const_431_2;
    wire const_432_0;
    wire const_433_0;
    wire const_434_0;
    wire const_435_0;
    wire const_436_0;
    wire const_437_0;
    wire[255:0] const_438_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_440_0;
    wire const_441_0;
    wire const_442_0;
    wire const_443_0;
    wire const_444_0;
    wire[255:0] const_445_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_447_0;
    wire const_448_0;
    wire const_449_0;
    wire const_450_0;
    wire const_451_0;
    wire[255:0] const_452_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_454_0;
    wire const_455_0;
    wire const_456_0;
    wire const_457_0;
    wire const_458_0;
    wire[255:0] const_459_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_461_0;
    wire const_462_0;
    wire const_463_0;
    wire const_464_0;
    wire const_465_0;
    wire[255:0] const_466_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_468_0;
    wire const_469_0;
    wire const_470_0;
    wire const_471_0;
    wire const_472_0;
    wire[255:0] const_473_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_475_0;
    wire const_476_0;
    wire const_477_0;
    wire const_478_0;
    wire const_479_0;
    wire[255:0] const_480_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_482_0;
    wire const_483_0;
    wire const_484_0;
    wire const_485_0;
    wire const_486_0;
    wire[255:0] const_487_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_489_0;
    wire const_490_0;
    wire const_491_0;
    wire const_492_0;
    wire const_493_0;
    wire[255:0] const_494_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_496_0;
    wire const_497_0;
    wire const_498_0;
    wire const_499_0;
    wire const_500_0;
    wire[255:0] const_501_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_503_0;
    wire const_504_0;
    wire const_505_0;
    wire const_506_0;
    wire const_507_0;
    wire[255:0] const_508_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_510_0;
    wire const_511_0;
    wire const_512_0;
    wire const_513_0;
    wire const_514_0;
    wire[255:0] const_515_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire[3:0] const_517_5;
    wire const_518_1;
    wire const_520_0;
    wire const_521_0;
    wire[254:0] const_522_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_523_0;
    wire const_524_0;
    wire const_525_0;
    wire const_526_0;
    wire const_527_0;
    wire const_528_0;
    wire const_529_0;
    wire[255:0] const_530_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_533_0;
    wire const_534_0;
    wire[254:0] const_535_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_536_0;
    wire const_537_0;
    wire const_538_0;
    wire const_539_0;
    wire const_540_0;
    wire const_541_0;
    wire const_542_0;
    wire[255:0] const_543_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_546_0;
    wire const_547_0;
    wire[254:0] const_548_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_549_0;
    wire const_550_0;
    wire const_551_0;
    wire const_552_0;
    wire const_553_0;
    wire const_554_0;
    wire const_555_0;
    wire[255:0] const_556_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_559_0;
    wire const_560_0;
    wire[254:0] const_561_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_562_0;
    wire const_563_0;
    wire const_564_0;
    wire const_565_0;
    wire const_566_0;
    wire const_567_0;
    wire const_568_0;
    wire[255:0] const_569_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire[3:0] const_571_0;
    wire const_572_0;
    wire[3:0] const_573_0;
    wire const_574_0;
    wire const_575_0;
    wire const_577_0;
    wire const_578_0;
    wire[254:0] const_579_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_580_0;
    wire const_581_0;
    wire const_582_0;
    wire const_584_0;
    wire const_585_0;
    wire[254:0] const_586_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_587_0;
    wire const_588_0;
    wire const_589_0;
    wire const_591_0;
    wire const_592_0;
    wire[254:0] const_593_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_594_0;
    wire const_595_0;
    wire const_596_0;
    wire const_598_0;
    wire const_599_0;
    wire[254:0] const_600_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_601_0;
    wire const_602_0;
    wire const_603_0;
    wire const_605_0;
    wire const_606_0;
    wire[254:0] const_607_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_608_0;
    wire const_609_0;
    wire const_610_0;
    wire const_612_0;
    wire const_613_0;
    wire[254:0] const_614_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_615_0;
    wire const_616_0;
    wire const_617_0;
    wire const_619_0;
    wire const_620_0;
    wire[254:0] const_621_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_622_0;
    wire const_623_0;
    wire const_624_0;
    wire const_626_0;
    wire const_627_0;
    wire[254:0] const_628_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_629_0;
    wire const_630_0;
    wire[3:0] const_631_6;
    wire const_632_1;
    wire const_633_0;
    wire const_635_0;
    wire const_636_0;
    wire[254:0] const_637_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_638_0;
    wire const_639_0;
    wire const_640_0;
    wire const_642_0;
    wire const_643_0;
    wire[254:0] const_644_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_645_0;
    wire const_646_0;
    wire const_647_0;
    wire const_649_0;
    wire const_650_0;
    wire[254:0] const_651_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_652_0;
    wire const_653_0;
    wire const_654_0;
    wire const_656_0;
    wire const_657_0;
    wire[254:0] const_658_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_659_0;
    wire const_660_0;
    wire const_661_0;
    wire const_663_0;
    wire const_664_0;
    wire[254:0] const_665_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_666_0;
    wire const_667_0;
    wire const_668_0;
    wire const_670_0;
    wire const_671_0;
    wire[254:0] const_672_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_673_0;
    wire const_674_0;
    wire const_675_0;
    wire const_677_0;
    wire const_678_0;
    wire[254:0] const_679_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_680_0;
    wire const_681_0;
    wire const_682_0;
    wire const_684_0;
    wire const_685_0;
    wire[254:0] const_686_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_687_0;
    wire const_688_0;
    wire[3:0] const_689_3;
    wire const_690_1;
    wire const_691_0;
    wire const_692_0;
    wire const_693_0;
    wire const_694_0;
    wire const_695_0;
    wire[255:0] const_696_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_698_0;
    wire const_699_0;
    wire const_700_0;
    wire const_701_0;
    wire const_702_0;
    wire[255:0] const_703_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_705_0;
    wire const_706_0;
    wire const_707_0;
    wire const_708_0;
    wire const_709_0;
    wire[255:0] const_710_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire const_712_0;
    wire const_713_0;
    wire const_714_0;
    wire const_715_0;
    wire const_716_0;
    wire[255:0] const_717_57896044618658097711785492504343953926634992332820282019728792003956564819967;
    wire[3:0] const_719_0;
    wire[3:0] const_720_0;
    wire const_721_0;
    wire const_722_0;
    wire const_723_0;
    wire const_724_0;
    wire const_725_0;
    wire const_726_0;
    wire const_727_0;
    wire const_728_0;
    wire const_729_0;
    wire const_730_0;
    wire const_731_0;
    wire const_732_0;
    wire const_733_0;
    wire const_734_0;
    wire const_735_0;
    wire const_736_0;
    wire const_737_0;
    wire const_738_0;
    wire const_739_0;
    wire const_740_0;
    wire const_741_0;
    wire const_742_0;
    wire const_743_0;
    wire const_744_1;
    wire const_745_0;
    wire[1:0] const_746_2;
    wire const_747_0;
    wire[1:0] const_748_3;
    wire const_749_0;
    wire[3:0] const_750_15;
    wire const_751_0;
    wire[2:0] const_752_4;
    wire[2:0] const_753_5;
    wire[2:0] const_754_6;
    wire[2:0] const_755_7;
    wire[3:0] const_756_15;
    wire const_757_0;
    wire[3:0] const_758_8;
    wire const_759_0;
    wire[2:0] const_760_6;
    wire[2:0] const_761_7;
    wire[3:0] const_762_15;
    wire const_763_0;
    wire const_764_0;
    wire const_765_0;
    wire[2:0] const_766_1;
    wire const_767_1;
    wire const_768_0;
    wire[3:0] const_769_1;
    wire[2:0] const_770_2;
    wire[1:0] const_771_2;
    wire const_772_0;
    wire[3:0] const_773_1;
    wire[2:0] const_774_3;
    wire[1:0] const_775_3;
    wire const_776_0;
    wire[2:0] const_777_1;
    wire const_778_0;
    wire const_779_0;
    wire const_780_0;
    wire const_781_0;
    wire const_782_0;
    wire const_783_0;
    wire[2:0] my_calculator_ctrl;
    wire[3:0] my_calculator_in_x;
    wire[3:0] my_calculator_in_y;
    wire[3:0] my_calculator_out_z;
    wire[24:0] tmp1;
    wire[25:0] tmp2;
    wire[26:0] tmp3;
    wire[25:0] tmp4;
    wire tmp6;
    wire tmp8;
    wire tmp9;
    wire tmp10;
    wire tmp20;
    wire tmp21;
    wire tmp22;
    wire tmp23;
    wire tmp24;
    wire[255:0] tmp25;
    wire[255:0] tmp26;
    wire[255:0] tmp27;
    wire[255:0] tmp28;
    wire[255:0] tmp29;
    wire[255:0] tmp30;
    wire[255:0] tmp31;
    wire[255:0] tmp32;
    wire[1:0] tmp33;
    wire[2:0] tmp34;
    wire tmp35;
    wire tmp36;
    wire tmp37;
    wire tmp38;
    wire tmp39;
    wire tmp40;
    wire tmp41;
    wire tmp42;
    wire tmp43;
    wire tmp44;
    wire tmp45;
    wire tmp46;
    wire tmp47;
    wire tmp48;
    wire tmp49;
    wire tmp50;
    wire tmp51;
    wire tmp52;
    wire tmp53;
    wire tmp54;
    wire[1:0] tmp55;
    wire[2:0] tmp56;
    wire tmp57;
    wire tmp58;
    wire tmp59;
    wire tmp60;
    wire tmp61;
    wire tmp62;
    wire tmp63;
    wire tmp64;
    wire tmp65;
    wire[2:0] tmp66;
    wire[3:0] tmp67;
    wire tmp68;
    wire tmp69;
    wire tmp70;
    wire tmp71;
    wire tmp72;
    wire tmp73;
    wire tmp74;
    wire tmp75;
    wire tmp76;
    wire tmp77;
    wire tmp78;
    wire tmp79;
    wire tmp80;
    wire tmp81;
    wire tmp82;
    wire tmp83;
    wire tmp84;
    wire tmp85;
    wire tmp86;
    wire tmp87;
    wire tmp88;
    wire tmp89;
    wire tmp90;
    wire tmp91;
    wire tmp92;
    wire tmp93;
    wire tmp94;
    wire tmp95;
    wire tmp96;
    wire tmp97;
    wire[2:0] tmp98;
    wire[3:0] tmp99;
    wire tmp100;
    wire[1:0] tmp101;
    wire[3:0] tmp102;
    wire tmp103;
    wire tmp104;
    wire[1:0] tmp105;
    wire[3:0] tmp106;
    wire tmp107;
    wire tmp108;
    wire[254:0] tmp109;
    wire[255:0] tmp110;
    wire tmp111;
    wire[254:0] tmp112;
    wire[255:0] tmp113;
    wire tmp114;
    wire[256:0] tmp115;
    wire tmp116;
    wire tmp117;
    wire tmp118;
    wire tmp119;
    wire tmp120;
    wire tmp121;
    wire tmp122;
    wire tmp123;
    wire tmp124;
    wire[254:0] tmp125;
    wire[255:0] tmp126;
    wire[256:0] tmp127;
    wire tmp128;
    wire tmp129;
    wire tmp130;
    wire tmp131;
    wire tmp132;
    wire tmp133;
    wire tmp134;
    wire tmp135;
    wire tmp136;
    wire tmp137;
    wire[254:0] tmp138;
    wire[255:0] tmp139;
    wire[256:0] tmp140;
    wire tmp141;
    wire tmp142;
    wire tmp143;
    wire tmp144;
    wire tmp145;
    wire tmp146;
    wire tmp147;
    wire tmp148;
    wire[254:0] tmp149;
    wire[255:0] tmp150;
    wire tmp151;
    wire[256:0] tmp152;
    wire tmp153;
    wire tmp154;
    wire tmp155;
    wire tmp156;
    wire tmp157;
    wire tmp158;
    wire tmp159;
    wire tmp160;
    wire tmp161;
    wire tmp162;
    wire[255:0] tmp163;
    wire[255:0] tmp164;
    wire tmp165;
    wire tmp166;
    wire tmp167;
    wire tmp168;
    wire tmp169;
    wire tmp170;
    wire tmp171;
    wire tmp172;
    wire tmp173;
    wire[254:0] tmp174;
    wire[255:0] tmp175;
    wire tmp176;
    wire[254:0] tmp177;
    wire[255:0] tmp178;
    wire tmp179;
    wire[256:0] tmp180;
    wire tmp181;
    wire tmp182;
    wire tmp183;
    wire tmp184;
    wire tmp185;
    wire tmp186;
    wire tmp187;
    wire tmp188;
    wire tmp189;
    wire[254:0] tmp190;
    wire[255:0] tmp191;
    wire[256:0] tmp192;
    wire tmp193;
    wire tmp194;
    wire tmp195;
    wire tmp196;
    wire tmp197;
    wire tmp198;
    wire tmp199;
    wire tmp200;
    wire tmp201;
    wire tmp202;
    wire[254:0] tmp203;
    wire[255:0] tmp204;
    wire[256:0] tmp205;
    wire tmp206;
    wire tmp207;
    wire tmp208;
    wire tmp209;
    wire tmp210;
    wire tmp211;
    wire tmp212;
    wire tmp213;
    wire[254:0] tmp214;
    wire[255:0] tmp215;
    wire tmp216;
    wire[256:0] tmp217;
    wire tmp218;
    wire tmp219;
    wire tmp220;
    wire tmp221;
    wire tmp222;
    wire tmp223;
    wire tmp224;
    wire tmp225;
    wire tmp226;
    wire tmp227;
    wire[255:0] tmp228;
    wire[255:0] tmp229;
    wire tmp230;
    wire tmp231;
    wire tmp232;
    wire tmp233;
    wire tmp234;
    wire tmp235;
    wire tmp236;
    wire tmp237;
    wire tmp238;
    wire[254:0] tmp239;
    wire[255:0] tmp240;
    wire tmp241;
    wire[254:0] tmp242;
    wire[255:0] tmp243;
    wire tmp244;
    wire[256:0] tmp245;
    wire tmp246;
    wire tmp247;
    wire tmp248;
    wire tmp249;
    wire tmp250;
    wire tmp251;
    wire tmp252;
    wire tmp253;
    wire tmp254;
    wire[254:0] tmp255;
    wire[255:0] tmp256;
    wire[256:0] tmp257;
    wire tmp258;
    wire tmp259;
    wire tmp260;
    wire tmp261;
    wire tmp262;
    wire tmp263;
    wire tmp264;
    wire tmp265;
    wire tmp266;
    wire tmp267;
    wire[254:0] tmp268;
    wire[255:0] tmp269;
    wire[256:0] tmp270;
    wire tmp271;
    wire tmp272;
    wire tmp273;
    wire tmp274;
    wire tmp275;
    wire tmp276;
    wire tmp277;
    wire tmp278;
    wire[254:0] tmp279;
    wire[255:0] tmp280;
    wire tmp281;
    wire[256:0] tmp282;
    wire tmp283;
    wire tmp284;
    wire tmp285;
    wire tmp286;
    wire tmp287;
    wire tmp288;
    wire tmp289;
    wire tmp290;
    wire tmp291;
    wire tmp292;
    wire[255:0] tmp293;
    wire[255:0] tmp294;
    wire tmp295;
    wire tmp296;
    wire tmp297;
    wire tmp298;
    wire tmp299;
    wire tmp300;
    wire tmp301;
    wire tmp302;
    wire tmp303;
    wire[254:0] tmp304;
    wire[255:0] tmp305;
    wire tmp306;
    wire[254:0] tmp307;
    wire[255:0] tmp308;
    wire tmp309;
    wire[256:0] tmp310;
    wire tmp311;
    wire tmp312;
    wire tmp313;
    wire tmp314;
    wire tmp315;
    wire tmp316;
    wire tmp317;
    wire tmp318;
    wire tmp319;
    wire[254:0] tmp320;
    wire[255:0] tmp321;
    wire[256:0] tmp322;
    wire tmp323;
    wire tmp324;
    wire tmp325;
    wire tmp326;
    wire tmp327;
    wire tmp328;
    wire tmp329;
    wire tmp330;
    wire tmp331;
    wire tmp332;
    wire[254:0] tmp333;
    wire[255:0] tmp334;
    wire[256:0] tmp335;
    wire tmp336;
    wire tmp337;
    wire tmp338;
    wire tmp339;
    wire tmp340;
    wire tmp341;
    wire tmp342;
    wire tmp343;
    wire[254:0] tmp344;
    wire[255:0] tmp345;
    wire tmp346;
    wire[256:0] tmp347;
    wire tmp348;
    wire tmp349;
    wire tmp350;
    wire tmp351;
    wire tmp352;
    wire tmp353;
    wire tmp354;
    wire tmp355;
    wire tmp356;
    wire tmp357;
    wire[255:0] tmp358;
    wire[255:0] tmp359;
    wire tmp360;
    wire tmp361;
    wire tmp362;
    wire tmp363;
    wire tmp364;
    wire tmp365;
    wire tmp366;
    wire tmp367;
    wire tmp368;
    wire tmp369;
    wire[3:0] tmp370;
    wire tmp371;
    wire tmp372;
    wire[3:0] tmp373;
    wire tmp374;
    wire tmp375;
    wire tmp376;
    wire tmp377;
    wire tmp378;
    wire tmp379;
    wire tmp380;
    wire tmp381;
    wire tmp382;
    wire tmp383;
    wire tmp384;
    wire tmp385;
    wire tmp386;
    wire tmp387;
    wire tmp388;
    wire tmp389;
    wire tmp390;
    wire tmp391;
    wire tmp392;
    wire tmp393;
    wire tmp394;
    wire tmp395;
    wire tmp396;
    wire tmp397;
    wire tmp398;
    wire tmp399;
    wire tmp400;
    wire tmp401;
    wire tmp402;
    wire tmp403;
    wire tmp404;
    wire tmp405;
    wire tmp406;
    wire tmp407;
    wire tmp408;
    wire tmp409;
    wire tmp410;
    wire tmp411;
    wire tmp412;
    wire tmp413;
    wire tmp414;
    wire tmp415;
    wire tmp416;
    wire tmp417;
    wire tmp418;
    wire tmp419;
    wire tmp420;
    wire tmp421;
    wire tmp422;
    wire tmp423;
    wire tmp424;
    wire tmp425;
    wire tmp426;
    wire tmp427;
    wire tmp428;
    wire tmp429;
    wire tmp430;
    wire tmp431;
    wire tmp432;
    wire tmp433;
    wire tmp434;
    wire tmp435;
    wire tmp436;
    wire tmp437;
    wire tmp438;
    wire tmp439;
    wire tmp440;
    wire tmp441;
    wire tmp442;
    wire tmp443;
    wire tmp444;
    wire tmp445;
    wire tmp446;
    wire tmp447;
    wire tmp448;
    wire tmp449;
    wire tmp450;
    wire tmp451;
    wire tmp452;
    wire tmp453;
    wire tmp454;
    wire tmp455;
    wire tmp456;
    wire tmp457;
    wire tmp458;
    wire tmp459;
    wire tmp460;
    wire tmp461;
    wire tmp462;
    wire tmp463;
    wire tmp464;
    wire[3:0] tmp465;
    wire tmp466;
    wire tmp467;
    wire[3:0] tmp468;
    wire tmp469;
    wire tmp470;
    wire tmp471;
    wire tmp472;
    wire[256:0] tmp473;
    wire tmp474;
    wire tmp475;
    wire[256:0] tmp476;
    wire[257:0] tmp477;
    wire[256:0] tmp478;
    wire[255:0] tmp479;
    wire tmp480;
    wire[254:0] tmp481;
    wire[255:0] tmp482;
    wire tmp483;
    wire[256:0] tmp484;
    wire tmp485;
    wire tmp486;
    wire tmp487;
    wire tmp488;
    wire tmp489;
    wire tmp490;
    wire tmp491;
    wire tmp492;
    wire[254:0] tmp493;
    wire[255:0] tmp494;
    wire tmp495;
    wire[256:0] tmp496;
    wire tmp497;
    wire tmp498;
    wire tmp499;
    wire tmp500;
    wire tmp501;
    wire tmp502;
    wire tmp503;
    wire tmp504;
    wire tmp505;
    wire tmp506;
    wire[254:0] tmp507;
    wire[255:0] tmp508;
    wire[256:0] tmp509;
    wire tmp510;
    wire tmp511;
    wire tmp512;
    wire tmp513;
    wire tmp514;
    wire tmp515;
    wire tmp516;
    wire tmp517;
    wire tmp518;
    wire tmp519;
    wire tmp520;
    wire tmp521;
    wire[254:0] tmp522;
    wire[255:0] tmp523;
    wire[256:0] tmp524;
    wire tmp525;
    wire tmp526;
    wire tmp527;
    wire tmp528;
    wire tmp529;
    wire tmp530;
    wire tmp531;
    wire tmp532;
    wire tmp533;
    wire[254:0] tmp534;
    wire[255:0] tmp535;
    wire[256:0] tmp536;
    wire tmp537;
    wire tmp538;
    wire tmp539;
    wire tmp540;
    wire tmp541;
    wire tmp542;
    wire tmp543;
    wire tmp544;
    wire tmp545;
    wire[254:0] tmp546;
    wire[255:0] tmp547;
    wire tmp548;
    wire[256:0] tmp549;
    wire tmp550;
    wire tmp551;
    wire tmp552;
    wire tmp553;
    wire tmp554;
    wire tmp555;
    wire tmp556;
    wire tmp557;
    wire tmp558;
    wire tmp559;
    wire[255:0] tmp560;
    wire[255:0] tmp561;
    wire tmp562;
    wire tmp563;
    wire tmp564;
    wire tmp565;
    wire tmp566;
    wire tmp567;
    wire tmp568;
    wire tmp569;
    wire tmp570;
    wire tmp571;
    wire tmp572;
    wire tmp573;
    wire tmp574;
    wire tmp575;
    wire tmp576;
    wire tmp577;
    wire tmp578;
    wire tmp579;
    wire tmp580;
    wire tmp581;
    wire tmp582;
    wire tmp583;
    wire tmp584;
    wire tmp585;
    wire tmp586;
    wire tmp587;
    wire tmp588;
    wire tmp589;
    wire[256:0] tmp590;
    wire tmp591;
    wire tmp592;
    wire[256:0] tmp593;
    wire[257:0] tmp594;
    wire[256:0] tmp595;
    wire[255:0] tmp596;
    wire tmp597;
    wire[254:0] tmp598;
    wire[255:0] tmp599;
    wire tmp600;
    wire[256:0] tmp601;
    wire tmp602;
    wire tmp603;
    wire tmp604;
    wire tmp605;
    wire tmp606;
    wire tmp607;
    wire tmp608;
    wire tmp609;
    wire[254:0] tmp610;
    wire[255:0] tmp611;
    wire tmp612;
    wire[256:0] tmp613;
    wire tmp614;
    wire tmp615;
    wire tmp616;
    wire tmp617;
    wire tmp618;
    wire tmp619;
    wire tmp620;
    wire tmp621;
    wire tmp622;
    wire tmp623;
    wire[254:0] tmp624;
    wire[255:0] tmp625;
    wire[256:0] tmp626;
    wire tmp627;
    wire tmp628;
    wire tmp629;
    wire tmp630;
    wire tmp631;
    wire tmp632;
    wire tmp633;
    wire tmp634;
    wire tmp635;
    wire tmp636;
    wire tmp637;
    wire tmp638;
    wire[254:0] tmp639;
    wire[255:0] tmp640;
    wire[256:0] tmp641;
    wire tmp642;
    wire tmp643;
    wire tmp644;
    wire tmp645;
    wire tmp646;
    wire tmp647;
    wire tmp648;
    wire tmp649;
    wire tmp650;
    wire[254:0] tmp651;
    wire[255:0] tmp652;
    wire[256:0] tmp653;
    wire tmp654;
    wire tmp655;
    wire tmp656;
    wire tmp657;
    wire tmp658;
    wire tmp659;
    wire tmp660;
    wire tmp661;
    wire tmp662;
    wire[254:0] tmp663;
    wire[255:0] tmp664;
    wire tmp665;
    wire[256:0] tmp666;
    wire tmp667;
    wire tmp668;
    wire tmp669;
    wire tmp670;
    wire tmp671;
    wire tmp672;
    wire tmp673;
    wire tmp674;
    wire tmp675;
    wire tmp676;
    wire[255:0] tmp677;
    wire[255:0] tmp678;
    wire tmp679;
    wire tmp680;
    wire tmp681;
    wire tmp682;
    wire tmp683;
    wire tmp684;
    wire tmp685;
    wire tmp686;
    wire tmp687;
    wire tmp688;
    wire tmp689;
    wire tmp690;
    wire tmp691;
    wire tmp692;
    wire tmp693;
    wire tmp694;
    wire tmp695;
    wire tmp696;
    wire tmp697;
    wire tmp698;
    wire tmp699;
    wire tmp700;
    wire tmp701;
    wire tmp702;
    wire tmp703;
    wire tmp704;
    wire tmp705;
    wire tmp706;
    wire[256:0] tmp707;
    wire tmp708;
    wire tmp709;
    wire[256:0] tmp710;
    wire[257:0] tmp711;
    wire[256:0] tmp712;
    wire[255:0] tmp713;
    wire tmp714;
    wire[254:0] tmp715;
    wire[255:0] tmp716;
    wire tmp717;
    wire[256:0] tmp718;
    wire tmp719;
    wire tmp720;
    wire tmp721;
    wire tmp722;
    wire tmp723;
    wire tmp724;
    wire tmp725;
    wire tmp726;
    wire[254:0] tmp727;
    wire[255:0] tmp728;
    wire tmp729;
    wire[256:0] tmp730;
    wire tmp731;
    wire tmp732;
    wire tmp733;
    wire tmp734;
    wire tmp735;
    wire tmp736;
    wire tmp737;
    wire tmp738;
    wire tmp739;
    wire tmp740;
    wire[254:0] tmp741;
    wire[255:0] tmp742;
    wire[256:0] tmp743;
    wire tmp744;
    wire tmp745;
    wire tmp746;
    wire tmp747;
    wire tmp748;
    wire tmp749;
    wire tmp750;
    wire tmp751;
    wire tmp752;
    wire tmp753;
    wire tmp754;
    wire tmp755;
    wire[254:0] tmp756;
    wire[255:0] tmp757;
    wire[256:0] tmp758;
    wire tmp759;
    wire tmp760;
    wire tmp761;
    wire tmp762;
    wire tmp763;
    wire tmp764;
    wire tmp765;
    wire tmp766;
    wire tmp767;
    wire[254:0] tmp768;
    wire[255:0] tmp769;
    wire[256:0] tmp770;
    wire tmp771;
    wire tmp772;
    wire tmp773;
    wire tmp774;
    wire tmp775;
    wire tmp776;
    wire tmp777;
    wire tmp778;
    wire tmp779;
    wire[254:0] tmp780;
    wire[255:0] tmp781;
    wire tmp782;
    wire[256:0] tmp783;
    wire tmp784;
    wire tmp785;
    wire tmp786;
    wire tmp787;
    wire tmp788;
    wire tmp789;
    wire tmp790;
    wire tmp791;
    wire tmp792;
    wire tmp793;
    wire[255:0] tmp794;
    wire[255:0] tmp795;
    wire tmp796;
    wire tmp797;
    wire tmp798;
    wire tmp799;
    wire tmp800;
    wire tmp801;
    wire tmp802;
    wire tmp803;
    wire tmp804;
    wire tmp805;
    wire tmp806;
    wire tmp807;
    wire tmp808;
    wire tmp809;
    wire tmp810;
    wire tmp811;
    wire tmp812;
    wire tmp813;
    wire tmp814;
    wire tmp815;
    wire tmp816;
    wire tmp817;
    wire tmp818;
    wire tmp819;
    wire tmp820;
    wire tmp821;
    wire tmp822;
    wire tmp823;
    wire[256:0] tmp824;
    wire tmp825;
    wire tmp826;
    wire[256:0] tmp827;
    wire[257:0] tmp828;
    wire[256:0] tmp829;
    wire[255:0] tmp830;
    wire tmp831;
    wire[254:0] tmp832;
    wire[255:0] tmp833;
    wire tmp834;
    wire[256:0] tmp835;
    wire tmp836;
    wire tmp837;
    wire tmp838;
    wire tmp839;
    wire tmp840;
    wire tmp841;
    wire tmp842;
    wire tmp843;
    wire[254:0] tmp844;
    wire[255:0] tmp845;
    wire tmp846;
    wire[256:0] tmp847;
    wire tmp848;
    wire tmp849;
    wire tmp850;
    wire tmp851;
    wire tmp852;
    wire tmp853;
    wire tmp854;
    wire tmp855;
    wire tmp856;
    wire tmp857;
    wire[254:0] tmp858;
    wire[255:0] tmp859;
    wire[256:0] tmp860;
    wire tmp861;
    wire tmp862;
    wire tmp863;
    wire tmp864;
    wire tmp865;
    wire tmp866;
    wire tmp867;
    wire tmp868;
    wire tmp869;
    wire tmp870;
    wire tmp871;
    wire tmp872;
    wire[254:0] tmp873;
    wire[255:0] tmp874;
    wire[256:0] tmp875;
    wire tmp876;
    wire tmp877;
    wire tmp878;
    wire tmp879;
    wire tmp880;
    wire tmp881;
    wire tmp882;
    wire tmp883;
    wire tmp884;
    wire[254:0] tmp885;
    wire[255:0] tmp886;
    wire[256:0] tmp887;
    wire tmp888;
    wire tmp889;
    wire tmp890;
    wire tmp891;
    wire tmp892;
    wire tmp893;
    wire tmp894;
    wire tmp895;
    wire tmp896;
    wire[254:0] tmp897;
    wire[255:0] tmp898;
    wire tmp899;
    wire[256:0] tmp900;
    wire tmp901;
    wire tmp902;
    wire tmp903;
    wire tmp904;
    wire tmp905;
    wire tmp906;
    wire tmp907;
    wire tmp908;
    wire tmp909;
    wire tmp910;
    wire[255:0] tmp911;
    wire[255:0] tmp912;
    wire tmp913;
    wire tmp914;
    wire tmp915;
    wire tmp916;
    wire tmp917;
    wire tmp918;
    wire tmp919;
    wire tmp920;
    wire tmp921;
    wire tmp922;
    wire tmp923;
    wire tmp924;
    wire tmp925;
    wire tmp926;
    wire tmp927;
    wire tmp928;
    wire tmp929;
    wire tmp930;
    wire tmp931;
    wire tmp932;
    wire tmp933;
    wire tmp934;
    wire tmp935;
    wire tmp936;
    wire tmp937;
    wire tmp938;
    wire tmp939;
    wire tmp940;
    wire[254:0] tmp941;
    wire[255:0] tmp942;
    wire[256:0] tmp943;
    wire[1:0] tmp944;
    wire[256:0] tmp945;
    wire[256:0] tmp946;
    wire[255:0] tmp947;
    wire tmp948;
    wire tmp949;
    wire tmp950;
    wire tmp951;
    wire tmp952;
    wire tmp953;
    wire tmp954;
    wire tmp955;
    wire tmp956;
    wire tmp957;
    wire tmp958;
    wire tmp959;
    wire tmp960;
    wire tmp961;
    wire tmp962;
    wire tmp963;
    wire[254:0] tmp964;
    wire[255:0] tmp965;
    wire[256:0] tmp966;
    wire[1:0] tmp967;
    wire[256:0] tmp968;
    wire[256:0] tmp969;
    wire[255:0] tmp970;
    wire tmp971;
    wire tmp972;
    wire tmp973;
    wire tmp974;
    wire tmp975;
    wire tmp976;
    wire tmp977;
    wire tmp978;
    wire tmp979;
    wire tmp980;
    wire tmp981;
    wire tmp982;
    wire tmp983;
    wire tmp984;
    wire tmp985;
    wire tmp986;
    wire[254:0] tmp987;
    wire[255:0] tmp988;
    wire[256:0] tmp989;
    wire[1:0] tmp990;
    wire[256:0] tmp991;
    wire[256:0] tmp992;
    wire[255:0] tmp993;
    wire tmp994;
    wire tmp995;
    wire tmp996;
    wire tmp997;
    wire tmp998;
    wire tmp999;
    wire tmp1000;
    wire tmp1001;
    wire tmp1002;
    wire tmp1003;
    wire tmp1004;
    wire tmp1005;
    wire tmp1006;
    wire tmp1007;
    wire tmp1008;
    wire tmp1009;
    wire[254:0] tmp1010;
    wire[255:0] tmp1011;
    wire[256:0] tmp1012;
    wire[1:0] tmp1013;
    wire[256:0] tmp1014;
    wire[256:0] tmp1015;
    wire[255:0] tmp1016;
    wire tmp1017;
    wire tmp1018;
    wire tmp1019;
    wire tmp1020;
    wire tmp1021;
    wire tmp1022;
    wire tmp1023;
    wire tmp1024;
    wire tmp1025;
    wire tmp1026;
    wire tmp1027;
    wire tmp1028;
    wire tmp1029;
    wire tmp1030;
    wire tmp1031;
    wire tmp1032;
    wire[2:0] tmp1033;
    wire tmp1034;
    wire tmp1035;
    wire tmp1036;
    wire tmp1037;
    wire tmp1038;
    wire tmp1039;
    wire tmp1040;
    wire tmp1041;
    wire tmp1042;
    wire tmp1043;
    wire tmp1044;
    wire tmp1045;
    wire tmp1046;
    wire[2:0] tmp1047;
    wire[3:0] tmp1048;
    wire tmp1049;
    wire tmp1050;
    wire tmp1051;
    wire tmp1052;
    wire tmp1053;
    wire tmp1054;
    wire tmp1055;
    wire tmp1056;
    wire tmp1057;
    wire tmp1058;
    wire tmp1059;
    wire tmp1060;
    wire tmp1061;
    wire tmp1062;
    wire tmp1063;
    wire tmp1064;
    wire tmp1065;
    wire tmp1066;
    wire tmp1067;
    wire tmp1068;
    wire tmp1069;
    wire tmp1070;
    wire tmp1071;
    wire tmp1072;
    wire tmp1073;
    wire tmp1074;
    wire tmp1075;
    wire tmp1076;
    wire tmp1077;
    wire tmp1078;
    wire tmp1079;
    wire tmp1080;
    wire tmp1081;
    wire tmp1082;
    wire tmp1083;
    wire tmp1084;
    wire tmp1085;
    wire tmp1086;
    wire[2:0] tmp1087;
    wire[3:0] tmp1088;
    wire tmp1089;
    wire[1:0] tmp1090;
    wire[3:0] tmp1091;
    wire tmp1092;
    wire tmp1093;
    wire[1:0] tmp1094;
    wire[3:0] tmp1095;
    wire tmp1096;
    wire tmp1097;
    wire[254:0] tmp1098;
    wire[255:0] tmp1099;
    wire tmp1100;
    wire[254:0] tmp1101;
    wire[255:0] tmp1102;
    wire tmp1103;
    wire[256:0] tmp1104;
    wire tmp1105;
    wire tmp1106;
    wire tmp1107;
    wire tmp1108;
    wire tmp1109;
    wire tmp1110;
    wire tmp1111;
    wire tmp1112;
    wire tmp1113;
    wire[254:0] tmp1114;
    wire[255:0] tmp1115;
    wire[256:0] tmp1116;
    wire tmp1117;
    wire tmp1118;
    wire tmp1119;
    wire tmp1120;
    wire tmp1121;
    wire tmp1122;
    wire tmp1123;
    wire tmp1124;
    wire tmp1125;
    wire tmp1126;
    wire[254:0] tmp1127;
    wire[255:0] tmp1128;
    wire[256:0] tmp1129;
    wire tmp1130;
    wire tmp1131;
    wire tmp1132;
    wire tmp1133;
    wire tmp1134;
    wire tmp1135;
    wire tmp1136;
    wire tmp1137;
    wire[254:0] tmp1138;
    wire[255:0] tmp1139;
    wire tmp1140;
    wire[256:0] tmp1141;
    wire tmp1142;
    wire tmp1143;
    wire tmp1144;
    wire tmp1145;
    wire tmp1146;
    wire tmp1147;
    wire tmp1148;
    wire tmp1149;
    wire tmp1150;
    wire tmp1151;
    wire[255:0] tmp1152;
    wire[255:0] tmp1153;
    wire tmp1154;
    wire tmp1155;
    wire tmp1156;
    wire tmp1157;
    wire tmp1158;
    wire tmp1159;
    wire tmp1160;
    wire tmp1161;
    wire tmp1162;
    wire tmp1163;
    wire tmp1164;
    wire[254:0] tmp1165;
    wire[255:0] tmp1166;
    wire tmp1167;
    wire[254:0] tmp1168;
    wire[255:0] tmp1169;
    wire tmp1170;
    wire[256:0] tmp1171;
    wire tmp1172;
    wire tmp1173;
    wire tmp1174;
    wire tmp1175;
    wire tmp1176;
    wire tmp1177;
    wire tmp1178;
    wire tmp1179;
    wire tmp1180;
    wire[254:0] tmp1181;
    wire[255:0] tmp1182;
    wire[256:0] tmp1183;
    wire tmp1184;
    wire tmp1185;
    wire tmp1186;
    wire tmp1187;
    wire tmp1188;
    wire tmp1189;
    wire tmp1190;
    wire tmp1191;
    wire tmp1192;
    wire tmp1193;
    wire[254:0] tmp1194;
    wire[255:0] tmp1195;
    wire[256:0] tmp1196;
    wire tmp1197;
    wire tmp1198;
    wire tmp1199;
    wire tmp1200;
    wire tmp1201;
    wire tmp1202;
    wire tmp1203;
    wire tmp1204;
    wire[254:0] tmp1205;
    wire[255:0] tmp1206;
    wire tmp1207;
    wire[256:0] tmp1208;
    wire tmp1209;
    wire tmp1210;
    wire tmp1211;
    wire tmp1212;
    wire tmp1213;
    wire tmp1214;
    wire tmp1215;
    wire tmp1216;
    wire tmp1217;
    wire tmp1218;
    wire[255:0] tmp1219;
    wire[255:0] tmp1220;
    wire tmp1221;
    wire tmp1222;
    wire tmp1223;
    wire tmp1224;
    wire tmp1225;
    wire tmp1226;
    wire tmp1227;
    wire tmp1228;
    wire tmp1229;
    wire tmp1230;
    wire tmp1231;
    wire[254:0] tmp1232;
    wire[255:0] tmp1233;
    wire tmp1234;
    wire[254:0] tmp1235;
    wire[255:0] tmp1236;
    wire tmp1237;
    wire[256:0] tmp1238;
    wire tmp1239;
    wire tmp1240;
    wire tmp1241;
    wire tmp1242;
    wire tmp1243;
    wire tmp1244;
    wire tmp1245;
    wire tmp1246;
    wire tmp1247;
    wire[254:0] tmp1248;
    wire[255:0] tmp1249;
    wire[256:0] tmp1250;
    wire tmp1251;
    wire tmp1252;
    wire tmp1253;
    wire tmp1254;
    wire tmp1255;
    wire tmp1256;
    wire tmp1257;
    wire tmp1258;
    wire tmp1259;
    wire tmp1260;
    wire[254:0] tmp1261;
    wire[255:0] tmp1262;
    wire[256:0] tmp1263;
    wire tmp1264;
    wire tmp1265;
    wire tmp1266;
    wire tmp1267;
    wire tmp1268;
    wire tmp1269;
    wire tmp1270;
    wire tmp1271;
    wire[254:0] tmp1272;
    wire[255:0] tmp1273;
    wire tmp1274;
    wire[256:0] tmp1275;
    wire tmp1276;
    wire tmp1277;
    wire tmp1278;
    wire tmp1279;
    wire tmp1280;
    wire tmp1281;
    wire tmp1282;
    wire tmp1283;
    wire tmp1284;
    wire tmp1285;
    wire[255:0] tmp1286;
    wire[255:0] tmp1287;
    wire tmp1288;
    wire tmp1289;
    wire tmp1290;
    wire tmp1291;
    wire tmp1292;
    wire tmp1293;
    wire tmp1294;
    wire tmp1295;
    wire tmp1296;
    wire tmp1297;
    wire tmp1298;
    wire[254:0] tmp1299;
    wire[255:0] tmp1300;
    wire tmp1301;
    wire[254:0] tmp1302;
    wire[255:0] tmp1303;
    wire tmp1304;
    wire[256:0] tmp1305;
    wire tmp1306;
    wire tmp1307;
    wire tmp1308;
    wire tmp1309;
    wire tmp1310;
    wire tmp1311;
    wire tmp1312;
    wire tmp1313;
    wire tmp1314;
    wire[254:0] tmp1315;
    wire[255:0] tmp1316;
    wire[256:0] tmp1317;
    wire tmp1318;
    wire tmp1319;
    wire tmp1320;
    wire tmp1321;
    wire tmp1322;
    wire tmp1323;
    wire tmp1324;
    wire tmp1325;
    wire tmp1326;
    wire tmp1327;
    wire[254:0] tmp1328;
    wire[255:0] tmp1329;
    wire[256:0] tmp1330;
    wire tmp1331;
    wire tmp1332;
    wire tmp1333;
    wire tmp1334;
    wire tmp1335;
    wire tmp1336;
    wire tmp1337;
    wire tmp1338;
    wire[254:0] tmp1339;
    wire[255:0] tmp1340;
    wire tmp1341;
    wire[256:0] tmp1342;
    wire tmp1343;
    wire tmp1344;
    wire tmp1345;
    wire tmp1346;
    wire tmp1347;
    wire tmp1348;
    wire tmp1349;
    wire tmp1350;
    wire tmp1351;
    wire tmp1352;
    wire[255:0] tmp1353;
    wire[255:0] tmp1354;
    wire tmp1355;
    wire tmp1356;
    wire tmp1357;
    wire tmp1358;
    wire tmp1359;
    wire tmp1360;
    wire tmp1361;
    wire tmp1362;
    wire tmp1363;
    wire tmp1364;
    wire tmp1365;
    wire tmp1366;
    wire[3:0] tmp1367;
    wire tmp1368;
    wire tmp1369;
    wire[3:0] tmp1370;
    wire tmp1371;
    wire tmp1372;
    wire tmp1373;
    wire tmp1374;
    wire tmp1375;
    wire tmp1376;
    wire tmp1377;
    wire tmp1378;
    wire tmp1379;
    wire tmp1380;
    wire tmp1381;
    wire tmp1382;
    wire tmp1383;
    wire tmp1384;
    wire tmp1385;
    wire tmp1386;
    wire tmp1387;
    wire tmp1388;
    wire tmp1389;
    wire tmp1390;
    wire tmp1391;
    wire tmp1392;
    wire tmp1393;
    wire tmp1394;
    wire tmp1395;
    wire tmp1396;
    wire tmp1397;
    wire tmp1398;
    wire tmp1399;
    wire tmp1400;
    wire tmp1401;
    wire tmp1402;
    wire tmp1403;
    wire tmp1404;
    wire tmp1405;
    wire tmp1406;
    wire tmp1407;
    wire tmp1408;
    wire tmp1409;
    wire tmp1410;
    wire tmp1411;
    wire tmp1412;
    wire tmp1413;
    wire tmp1414;
    wire tmp1415;
    wire tmp1416;
    wire tmp1417;
    wire tmp1418;
    wire tmp1419;
    wire tmp1420;
    wire tmp1421;
    wire tmp1422;
    wire tmp1423;
    wire tmp1424;
    wire tmp1425;
    wire tmp1426;
    wire tmp1427;
    wire tmp1428;
    wire tmp1429;
    wire tmp1430;
    wire tmp1431;
    wire tmp1432;
    wire tmp1433;
    wire tmp1434;
    wire tmp1435;
    wire tmp1436;
    wire tmp1437;
    wire tmp1438;
    wire tmp1439;
    wire tmp1440;
    wire tmp1441;
    wire tmp1442;
    wire tmp1443;
    wire tmp1444;
    wire tmp1445;
    wire tmp1446;
    wire tmp1447;
    wire tmp1448;
    wire tmp1449;
    wire tmp1450;
    wire tmp1451;
    wire tmp1452;
    wire tmp1453;
    wire tmp1454;
    wire tmp1455;
    wire tmp1456;
    wire tmp1457;
    wire tmp1458;
    wire tmp1459;
    wire tmp1460;
    wire tmp1461;
    wire tmp1462;
    wire tmp1463;
    wire tmp1464;
    wire tmp1465;
    wire tmp1466;
    wire tmp1467;
    wire tmp1468;
    wire tmp1469;
    wire tmp1470;
    wire tmp1471;
    wire tmp1472;
    wire tmp1473;
    wire tmp1474;
    wire tmp1475;
    wire tmp1476;
    wire tmp1477;
    wire[3:0] tmp1478;
    wire tmp1479;
    wire tmp1480;
    wire[3:0] tmp1481;
    wire tmp1482;
    wire tmp1483;
    wire tmp1484;
    wire tmp1485;
    wire[256:0] tmp1486;
    wire tmp1487;
    wire tmp1488;
    wire[256:0] tmp1489;
    wire[257:0] tmp1490;
    wire[256:0] tmp1491;
    wire[255:0] tmp1492;
    wire tmp1493;
    wire[254:0] tmp1494;
    wire[255:0] tmp1495;
    wire tmp1496;
    wire[256:0] tmp1497;
    wire tmp1498;
    wire tmp1499;
    wire tmp1500;
    wire tmp1501;
    wire tmp1502;
    wire tmp1503;
    wire tmp1504;
    wire tmp1505;
    wire[254:0] tmp1506;
    wire[255:0] tmp1507;
    wire tmp1508;
    wire[256:0] tmp1509;
    wire tmp1510;
    wire tmp1511;
    wire tmp1512;
    wire tmp1513;
    wire tmp1514;
    wire tmp1515;
    wire tmp1516;
    wire tmp1517;
    wire tmp1518;
    wire tmp1519;
    wire[254:0] tmp1520;
    wire[255:0] tmp1521;
    wire[256:0] tmp1522;
    wire tmp1523;
    wire tmp1524;
    wire tmp1525;
    wire tmp1526;
    wire tmp1527;
    wire tmp1528;
    wire tmp1529;
    wire tmp1530;
    wire tmp1531;
    wire tmp1532;
    wire tmp1533;
    wire tmp1534;
    wire[254:0] tmp1535;
    wire[255:0] tmp1536;
    wire[256:0] tmp1537;
    wire tmp1538;
    wire tmp1539;
    wire tmp1540;
    wire tmp1541;
    wire tmp1542;
    wire tmp1543;
    wire tmp1544;
    wire tmp1545;
    wire tmp1546;
    wire[254:0] tmp1547;
    wire[255:0] tmp1548;
    wire[256:0] tmp1549;
    wire tmp1550;
    wire tmp1551;
    wire tmp1552;
    wire tmp1553;
    wire tmp1554;
    wire tmp1555;
    wire tmp1556;
    wire tmp1557;
    wire tmp1558;
    wire[254:0] tmp1559;
    wire[255:0] tmp1560;
    wire tmp1561;
    wire[256:0] tmp1562;
    wire tmp1563;
    wire tmp1564;
    wire tmp1565;
    wire tmp1566;
    wire tmp1567;
    wire tmp1568;
    wire tmp1569;
    wire tmp1570;
    wire tmp1571;
    wire tmp1572;
    wire[255:0] tmp1573;
    wire[255:0] tmp1574;
    wire tmp1575;
    wire tmp1576;
    wire tmp1577;
    wire tmp1578;
    wire tmp1579;
    wire tmp1580;
    wire tmp1581;
    wire tmp1582;
    wire tmp1583;
    wire tmp1584;
    wire tmp1585;
    wire tmp1586;
    wire tmp1587;
    wire tmp1588;
    wire tmp1589;
    wire tmp1590;
    wire tmp1591;
    wire tmp1592;
    wire tmp1593;
    wire tmp1594;
    wire tmp1595;
    wire tmp1596;
    wire tmp1597;
    wire tmp1598;
    wire tmp1599;
    wire tmp1600;
    wire tmp1601;
    wire tmp1602;
    wire tmp1603;
    wire tmp1604;
    wire tmp1605;
    wire tmp1606;
    wire[256:0] tmp1607;
    wire tmp1608;
    wire tmp1609;
    wire[256:0] tmp1610;
    wire[257:0] tmp1611;
    wire[256:0] tmp1612;
    wire[255:0] tmp1613;
    wire tmp1614;
    wire[254:0] tmp1615;
    wire[255:0] tmp1616;
    wire tmp1617;
    wire[256:0] tmp1618;
    wire tmp1619;
    wire tmp1620;
    wire tmp1621;
    wire tmp1622;
    wire tmp1623;
    wire tmp1624;
    wire tmp1625;
    wire tmp1626;
    wire[254:0] tmp1627;
    wire[255:0] tmp1628;
    wire tmp1629;
    wire[256:0] tmp1630;
    wire tmp1631;
    wire tmp1632;
    wire tmp1633;
    wire tmp1634;
    wire tmp1635;
    wire tmp1636;
    wire tmp1637;
    wire tmp1638;
    wire tmp1639;
    wire tmp1640;
    wire[254:0] tmp1641;
    wire[255:0] tmp1642;
    wire[256:0] tmp1643;
    wire tmp1644;
    wire tmp1645;
    wire tmp1646;
    wire tmp1647;
    wire tmp1648;
    wire tmp1649;
    wire tmp1650;
    wire tmp1651;
    wire tmp1652;
    wire tmp1653;
    wire tmp1654;
    wire tmp1655;
    wire[254:0] tmp1656;
    wire[255:0] tmp1657;
    wire[256:0] tmp1658;
    wire tmp1659;
    wire tmp1660;
    wire tmp1661;
    wire tmp1662;
    wire tmp1663;
    wire tmp1664;
    wire tmp1665;
    wire tmp1666;
    wire tmp1667;
    wire[254:0] tmp1668;
    wire[255:0] tmp1669;
    wire[256:0] tmp1670;
    wire tmp1671;
    wire tmp1672;
    wire tmp1673;
    wire tmp1674;
    wire tmp1675;
    wire tmp1676;
    wire tmp1677;
    wire tmp1678;
    wire tmp1679;
    wire[254:0] tmp1680;
    wire[255:0] tmp1681;
    wire tmp1682;
    wire[256:0] tmp1683;
    wire tmp1684;
    wire tmp1685;
    wire tmp1686;
    wire tmp1687;
    wire tmp1688;
    wire tmp1689;
    wire tmp1690;
    wire tmp1691;
    wire tmp1692;
    wire tmp1693;
    wire[255:0] tmp1694;
    wire[255:0] tmp1695;
    wire tmp1696;
    wire tmp1697;
    wire tmp1698;
    wire tmp1699;
    wire tmp1700;
    wire tmp1701;
    wire tmp1702;
    wire tmp1703;
    wire tmp1704;
    wire tmp1705;
    wire tmp1706;
    wire tmp1707;
    wire tmp1708;
    wire tmp1709;
    wire tmp1710;
    wire tmp1711;
    wire tmp1712;
    wire tmp1713;
    wire tmp1714;
    wire tmp1715;
    wire tmp1716;
    wire tmp1717;
    wire tmp1718;
    wire tmp1719;
    wire tmp1720;
    wire tmp1721;
    wire tmp1722;
    wire tmp1723;
    wire tmp1724;
    wire tmp1725;
    wire tmp1726;
    wire tmp1727;
    wire[256:0] tmp1728;
    wire tmp1729;
    wire tmp1730;
    wire[256:0] tmp1731;
    wire[257:0] tmp1732;
    wire[256:0] tmp1733;
    wire[255:0] tmp1734;
    wire tmp1735;
    wire[254:0] tmp1736;
    wire[255:0] tmp1737;
    wire tmp1738;
    wire[256:0] tmp1739;
    wire tmp1740;
    wire tmp1741;
    wire tmp1742;
    wire tmp1743;
    wire tmp1744;
    wire tmp1745;
    wire tmp1746;
    wire tmp1747;
    wire[254:0] tmp1748;
    wire[255:0] tmp1749;
    wire tmp1750;
    wire[256:0] tmp1751;
    wire tmp1752;
    wire tmp1753;
    wire tmp1754;
    wire tmp1755;
    wire tmp1756;
    wire tmp1757;
    wire tmp1758;
    wire tmp1759;
    wire tmp1760;
    wire tmp1761;
    wire[254:0] tmp1762;
    wire[255:0] tmp1763;
    wire[256:0] tmp1764;
    wire tmp1765;
    wire tmp1766;
    wire tmp1767;
    wire tmp1768;
    wire tmp1769;
    wire tmp1770;
    wire tmp1771;
    wire tmp1772;
    wire tmp1773;
    wire tmp1774;
    wire tmp1775;
    wire tmp1776;
    wire[254:0] tmp1777;
    wire[255:0] tmp1778;
    wire[256:0] tmp1779;
    wire tmp1780;
    wire tmp1781;
    wire tmp1782;
    wire tmp1783;
    wire tmp1784;
    wire tmp1785;
    wire tmp1786;
    wire tmp1787;
    wire tmp1788;
    wire[254:0] tmp1789;
    wire[255:0] tmp1790;
    wire[256:0] tmp1791;
    wire tmp1792;
    wire tmp1793;
    wire tmp1794;
    wire tmp1795;
    wire tmp1796;
    wire tmp1797;
    wire tmp1798;
    wire tmp1799;
    wire tmp1800;
    wire[254:0] tmp1801;
    wire[255:0] tmp1802;
    wire tmp1803;
    wire[256:0] tmp1804;
    wire tmp1805;
    wire tmp1806;
    wire tmp1807;
    wire tmp1808;
    wire tmp1809;
    wire tmp1810;
    wire tmp1811;
    wire tmp1812;
    wire tmp1813;
    wire tmp1814;
    wire[255:0] tmp1815;
    wire[255:0] tmp1816;
    wire tmp1817;
    wire tmp1818;
    wire tmp1819;
    wire tmp1820;
    wire tmp1821;
    wire tmp1822;
    wire tmp1823;
    wire tmp1824;
    wire tmp1825;
    wire tmp1826;
    wire tmp1827;
    wire tmp1828;
    wire tmp1829;
    wire tmp1830;
    wire tmp1831;
    wire tmp1832;
    wire tmp1833;
    wire tmp1834;
    wire tmp1835;
    wire tmp1836;
    wire tmp1837;
    wire tmp1838;
    wire tmp1839;
    wire tmp1840;
    wire tmp1841;
    wire tmp1842;
    wire tmp1843;
    wire tmp1844;
    wire tmp1845;
    wire tmp1846;
    wire tmp1847;
    wire tmp1848;
    wire[256:0] tmp1849;
    wire tmp1850;
    wire tmp1851;
    wire[256:0] tmp1852;
    wire[257:0] tmp1853;
    wire[256:0] tmp1854;
    wire[255:0] tmp1855;
    wire tmp1856;
    wire[254:0] tmp1857;
    wire[255:0] tmp1858;
    wire tmp1859;
    wire[256:0] tmp1860;
    wire tmp1861;
    wire tmp1862;
    wire tmp1863;
    wire tmp1864;
    wire tmp1865;
    wire tmp1866;
    wire tmp1867;
    wire tmp1868;
    wire[254:0] tmp1869;
    wire[255:0] tmp1870;
    wire tmp1871;
    wire[256:0] tmp1872;
    wire tmp1873;
    wire tmp1874;
    wire tmp1875;
    wire tmp1876;
    wire tmp1877;
    wire tmp1878;
    wire tmp1879;
    wire tmp1880;
    wire tmp1881;
    wire tmp1882;
    wire[254:0] tmp1883;
    wire[255:0] tmp1884;
    wire[256:0] tmp1885;
    wire tmp1886;
    wire tmp1887;
    wire tmp1888;
    wire tmp1889;
    wire tmp1890;
    wire tmp1891;
    wire tmp1892;
    wire tmp1893;
    wire tmp1894;
    wire tmp1895;
    wire tmp1896;
    wire tmp1897;
    wire[254:0] tmp1898;
    wire[255:0] tmp1899;
    wire[256:0] tmp1900;
    wire tmp1901;
    wire tmp1902;
    wire tmp1903;
    wire tmp1904;
    wire tmp1905;
    wire tmp1906;
    wire tmp1907;
    wire tmp1908;
    wire tmp1909;
    wire[254:0] tmp1910;
    wire[255:0] tmp1911;
    wire[256:0] tmp1912;
    wire tmp1913;
    wire tmp1914;
    wire tmp1915;
    wire tmp1916;
    wire tmp1917;
    wire tmp1918;
    wire tmp1919;
    wire tmp1920;
    wire tmp1921;
    wire[254:0] tmp1922;
    wire[255:0] tmp1923;
    wire tmp1924;
    wire[256:0] tmp1925;
    wire tmp1926;
    wire tmp1927;
    wire tmp1928;
    wire tmp1929;
    wire tmp1930;
    wire tmp1931;
    wire tmp1932;
    wire tmp1933;
    wire tmp1934;
    wire tmp1935;
    wire[255:0] tmp1936;
    wire[255:0] tmp1937;
    wire tmp1938;
    wire tmp1939;
    wire tmp1940;
    wire tmp1941;
    wire tmp1942;
    wire tmp1943;
    wire tmp1944;
    wire tmp1945;
    wire tmp1946;
    wire tmp1947;
    wire tmp1948;
    wire tmp1949;
    wire tmp1950;
    wire tmp1951;
    wire tmp1952;
    wire tmp1953;
    wire tmp1954;
    wire tmp1955;
    wire tmp1956;
    wire tmp1957;
    wire tmp1958;
    wire tmp1959;
    wire tmp1960;
    wire tmp1961;
    wire tmp1962;
    wire tmp1963;
    wire tmp1964;
    wire tmp1965;
    wire tmp1966;
    wire tmp1967;
    wire tmp1968;
    wire tmp1969;
    wire[254:0] tmp1970;
    wire[255:0] tmp1971;
    wire[256:0] tmp1972;
    wire[1:0] tmp1973;
    wire[256:0] tmp1974;
    wire[256:0] tmp1975;
    wire[255:0] tmp1976;
    wire tmp1977;
    wire tmp1978;
    wire tmp1979;
    wire tmp1980;
    wire tmp1981;
    wire tmp1982;
    wire tmp1983;
    wire tmp1984;
    wire tmp1985;
    wire tmp1986;
    wire tmp1987;
    wire tmp1988;
    wire tmp1989;
    wire tmp1990;
    wire tmp1991;
    wire tmp1992;
    wire tmp1993;
    wire tmp1994;
    wire[254:0] tmp1995;
    wire[255:0] tmp1996;
    wire[256:0] tmp1997;
    wire[1:0] tmp1998;
    wire[256:0] tmp1999;
    wire[256:0] tmp2000;
    wire[255:0] tmp2001;
    wire tmp2002;
    wire tmp2003;
    wire tmp2004;
    wire tmp2005;
    wire tmp2006;
    wire tmp2007;
    wire tmp2008;
    wire tmp2009;
    wire tmp2010;
    wire tmp2011;
    wire tmp2012;
    wire tmp2013;
    wire tmp2014;
    wire tmp2015;
    wire tmp2016;
    wire tmp2017;
    wire tmp2018;
    wire tmp2019;
    wire[254:0] tmp2020;
    wire[255:0] tmp2021;
    wire[256:0] tmp2022;
    wire[1:0] tmp2023;
    wire[256:0] tmp2024;
    wire[256:0] tmp2025;
    wire[255:0] tmp2026;
    wire tmp2027;
    wire tmp2028;
    wire tmp2029;
    wire tmp2030;
    wire tmp2031;
    wire tmp2032;
    wire tmp2033;
    wire tmp2034;
    wire tmp2035;
    wire tmp2036;
    wire tmp2037;
    wire tmp2038;
    wire tmp2039;
    wire tmp2040;
    wire tmp2041;
    wire tmp2042;
    wire tmp2043;
    wire tmp2044;
    wire[254:0] tmp2045;
    wire[255:0] tmp2046;
    wire[256:0] tmp2047;
    wire[1:0] tmp2048;
    wire[256:0] tmp2049;
    wire[256:0] tmp2050;
    wire[255:0] tmp2051;
    wire tmp2052;
    wire tmp2053;
    wire tmp2054;
    wire tmp2055;
    wire tmp2056;
    wire tmp2057;
    wire tmp2058;
    wire tmp2059;
    wire tmp2060;
    wire tmp2061;
    wire tmp2062;
    wire tmp2063;
    wire tmp2064;
    wire tmp2065;
    wire tmp2066;
    wire tmp2067;
    wire tmp2068;
    wire tmp2069;
    wire[2:0] tmp2070;
    wire tmp2071;
    wire tmp2072;
    wire tmp2073;
    wire[254:0] tmp2074;
    wire[255:0] tmp2075;
    wire[256:0] tmp2076;
    wire tmp2077;
    wire tmp2078;
    wire tmp2079;
    wire tmp2080;
    wire tmp2081;
    wire tmp2082;
    wire tmp2083;
    wire tmp2084;
    wire tmp2085;
    wire[254:0] tmp2086;
    wire[255:0] tmp2087;
    wire[256:0] tmp2088;
    wire tmp2089;
    wire tmp2090;
    wire tmp2091;
    wire tmp2092;
    wire tmp2093;
    wire tmp2094;
    wire tmp2095;
    wire tmp2096;
    wire tmp2097;
    wire tmp2098;
    wire[254:0] tmp2099;
    wire[255:0] tmp2100;
    wire[256:0] tmp2101;
    wire tmp2102;
    wire tmp2103;
    wire tmp2104;
    wire tmp2105;
    wire tmp2106;
    wire tmp2107;
    wire tmp2108;
    wire tmp2109;
    wire tmp2110;
    wire[254:0] tmp2111;
    wire[255:0] tmp2112;
    wire[256:0] tmp2113;
    wire tmp2114;
    wire tmp2115;
    wire tmp2116;
    wire tmp2117;
    wire tmp2118;
    wire tmp2119;
    wire tmp2120;
    wire tmp2121;
    wire tmp2122;
    wire tmp2123;
    wire tmp2124;
    wire[254:0] tmp2125;
    wire[255:0] tmp2126;
    wire[256:0] tmp2127;
    wire tmp2128;
    wire tmp2129;
    wire tmp2130;
    wire tmp2131;
    wire tmp2132;
    wire tmp2133;
    wire tmp2134;
    wire tmp2135;
    wire tmp2136;
    wire[254:0] tmp2137;
    wire[255:0] tmp2138;
    wire[256:0] tmp2139;
    wire tmp2140;
    wire tmp2141;
    wire tmp2142;
    wire tmp2143;
    wire tmp2144;
    wire tmp2145;
    wire tmp2146;
    wire tmp2147;
    wire tmp2148;
    wire tmp2149;
    wire tmp2150;
    wire tmp2151;
    wire tmp2152;
    wire tmp2153;
    wire tmp2154;
    wire tmp2155;
    wire tmp2156;
    wire tmp2157;
    wire tmp2158;
    wire[254:0] tmp2159;
    wire[255:0] tmp2160;
    wire[256:0] tmp2161;
    wire tmp2162;
    wire tmp2163;
    wire tmp2164;
    wire tmp2165;
    wire tmp2166;
    wire tmp2167;
    wire tmp2168;
    wire tmp2169;
    wire tmp2170;
    wire[254:0] tmp2171;
    wire[255:0] tmp2172;
    wire[256:0] tmp2173;
    wire tmp2174;
    wire tmp2175;
    wire tmp2176;
    wire tmp2177;
    wire tmp2178;
    wire tmp2179;
    wire tmp2180;
    wire tmp2181;
    wire tmp2182;
    wire tmp2183;
    wire[254:0] tmp2184;
    wire[255:0] tmp2185;
    wire[256:0] tmp2186;
    wire tmp2187;
    wire tmp2188;
    wire tmp2189;
    wire tmp2190;
    wire tmp2191;
    wire tmp2192;
    wire tmp2193;
    wire tmp2194;
    wire tmp2195;
    wire[254:0] tmp2196;
    wire[255:0] tmp2197;
    wire[256:0] tmp2198;
    wire tmp2199;
    wire tmp2200;
    wire tmp2201;
    wire tmp2202;
    wire tmp2203;
    wire tmp2204;
    wire tmp2205;
    wire tmp2206;
    wire tmp2207;
    wire tmp2208;
    wire tmp2209;
    wire[254:0] tmp2210;
    wire[255:0] tmp2211;
    wire[256:0] tmp2212;
    wire tmp2213;
    wire tmp2214;
    wire tmp2215;
    wire tmp2216;
    wire tmp2217;
    wire tmp2218;
    wire tmp2219;
    wire tmp2220;
    wire tmp2221;
    wire[254:0] tmp2222;
    wire[255:0] tmp2223;
    wire[256:0] tmp2224;
    wire tmp2225;
    wire tmp2226;
    wire tmp2227;
    wire tmp2228;
    wire tmp2229;
    wire tmp2230;
    wire tmp2231;
    wire tmp2232;
    wire tmp2233;
    wire tmp2234;
    wire tmp2235;
    wire tmp2236;
    wire tmp2237;
    wire tmp2238;
    wire tmp2239;
    wire tmp2240;
    wire tmp2241;
    wire[254:0] tmp2242;
    wire[255:0] tmp2243;
    wire tmp2244;
    wire[254:0] tmp2245;
    wire[255:0] tmp2246;
    wire tmp2247;
    wire tmp2248;
    wire[254:0] tmp2249;
    wire[255:0] tmp2250;
    wire tmp2251;
    wire tmp2252;
    wire[254:0] tmp2253;
    wire[255:0] tmp2254;
    wire tmp2255;
    wire tmp2256;
    wire tmp2257;
    wire tmp2258;
    wire tmp2259;
    wire tmp2260;
    wire tmp2261;
    wire tmp2262;
    wire tmp2263;
    wire tmp2264;
    wire tmp2265;
    wire tmp2266;
    wire tmp2267;
    wire tmp2268;
    wire tmp2269;
    wire tmp2270;
    wire tmp2271;
    wire tmp2272;
    wire tmp2273;
    wire tmp2274;
    wire tmp2275;
    wire tmp2276;
    wire tmp2277;
    wire tmp2278;
    wire tmp2279;
    wire tmp2280;
    wire tmp2281;
    wire tmp2282;
    wire tmp2283;
    wire tmp2284;
    wire tmp2285;
    wire tmp2286;
    wire tmp2287;
    wire tmp2288;
    wire tmp2289;
    wire tmp2290;
    wire tmp2291;
    wire tmp2292;
    wire tmp2293;
    wire[254:0] tmp2294;
    wire[255:0] tmp2295;
    wire[256:0] tmp2296;
    wire tmp2297;
    wire tmp2298;
    wire tmp2299;
    wire tmp2300;
    wire tmp2301;
    wire tmp2302;
    wire tmp2303;
    wire tmp2304;
    wire tmp2305;
    wire tmp2306;
    wire[254:0] tmp2307;
    wire[255:0] tmp2308;
    wire[256:0] tmp2309;
    wire tmp2310;
    wire tmp2311;
    wire tmp2312;
    wire tmp2313;
    wire tmp2314;
    wire tmp2315;
    wire tmp2316;
    wire tmp2317;
    wire tmp2318;
    wire[254:0] tmp2319;
    wire[255:0] tmp2320;
    wire[256:0] tmp2321;
    wire[1:0] tmp2322;
    wire[256:0] tmp2323;
    wire[256:0] tmp2324;
    wire[255:0] tmp2325;
    wire tmp2326;
    wire tmp2327;
    wire tmp2328;
    wire tmp2329;
    wire tmp2330;
    wire tmp2331;
    wire tmp2332;
    wire tmp2333;
    wire tmp2334;
    wire tmp2335;
    wire[254:0] tmp2336;
    wire[255:0] tmp2337;
    wire[256:0] tmp2338;
    wire[1:0] tmp2339;
    wire[256:0] tmp2340;
    wire[256:0] tmp2341;
    wire[255:0] tmp2342;
    wire tmp2343;
    wire tmp2344;
    wire tmp2345;
    wire tmp2346;
    wire tmp2347;
    wire tmp2348;
    wire tmp2349;
    wire tmp2350;
    wire tmp2351;
    wire tmp2352;
    wire[254:0] tmp2353;
    wire[255:0] tmp2354;
    wire[256:0] tmp2355;
    wire[1:0] tmp2356;
    wire[256:0] tmp2357;
    wire[256:0] tmp2358;
    wire[255:0] tmp2359;
    wire tmp2360;
    wire tmp2361;
    wire tmp2362;
    wire tmp2363;
    wire tmp2364;
    wire tmp2365;
    wire tmp2366;
    wire tmp2367;
    wire tmp2368;
    wire tmp2369;
    wire[254:0] tmp2370;
    wire[255:0] tmp2371;
    wire[256:0] tmp2372;
    wire[1:0] tmp2373;
    wire[256:0] tmp2374;
    wire[256:0] tmp2375;
    wire[255:0] tmp2376;
    wire tmp2377;
    wire tmp2378;
    wire tmp2379;
    wire tmp2380;
    wire tmp2381;
    wire tmp2382;
    wire tmp2383;
    wire tmp2384;
    wire tmp2385;
    wire tmp2386;
    wire[254:0] tmp2387;
    wire[255:0] tmp2388;
    wire[256:0] tmp2389;
    wire[1:0] tmp2390;
    wire[256:0] tmp2391;
    wire[256:0] tmp2392;
    wire[255:0] tmp2393;
    wire tmp2394;
    wire tmp2395;
    wire tmp2396;
    wire tmp2397;
    wire tmp2398;
    wire tmp2399;
    wire tmp2400;
    wire tmp2401;
    wire tmp2402;
    wire tmp2403;
    wire[254:0] tmp2404;
    wire[255:0] tmp2405;
    wire[256:0] tmp2406;
    wire[1:0] tmp2407;
    wire[256:0] tmp2408;
    wire[256:0] tmp2409;
    wire[255:0] tmp2410;
    wire tmp2411;
    wire tmp2412;
    wire tmp2413;
    wire tmp2414;
    wire tmp2415;
    wire tmp2416;
    wire tmp2417;
    wire tmp2418;
    wire tmp2419;
    wire tmp2420;
    wire[254:0] tmp2421;
    wire[255:0] tmp2422;
    wire[256:0] tmp2423;
    wire[1:0] tmp2424;
    wire[256:0] tmp2425;
    wire[256:0] tmp2426;
    wire[255:0] tmp2427;
    wire tmp2428;
    wire tmp2429;
    wire tmp2430;
    wire tmp2431;
    wire tmp2432;
    wire tmp2433;
    wire tmp2434;
    wire tmp2435;
    wire tmp2436;
    wire tmp2437;
    wire[254:0] tmp2438;
    wire[255:0] tmp2439;
    wire[256:0] tmp2440;
    wire[1:0] tmp2441;
    wire[256:0] tmp2442;
    wire[256:0] tmp2443;
    wire[255:0] tmp2444;
    wire tmp2445;
    wire tmp2446;
    wire tmp2447;
    wire tmp2448;
    wire tmp2449;
    wire tmp2450;
    wire tmp2451;
    wire tmp2452;
    wire tmp2453;
    wire tmp2454;
    wire tmp2455;
    wire[254:0] tmp2456;
    wire[255:0] tmp2457;
    wire[256:0] tmp2458;
    wire tmp2459;
    wire tmp2460;
    wire tmp2461;
    wire tmp2462;
    wire tmp2463;
    wire tmp2464;
    wire tmp2465;
    wire tmp2466;
    wire tmp2467;
    wire[254:0] tmp2468;
    wire[255:0] tmp2469;
    wire[256:0] tmp2470;
    wire tmp2471;
    wire tmp2472;
    wire tmp2473;
    wire tmp2474;
    wire tmp2475;
    wire tmp2476;
    wire tmp2477;
    wire tmp2478;
    wire tmp2479;
    wire tmp2480;
    wire tmp2481;
    wire tmp2482;
    wire tmp2483;
    wire tmp2484;
    wire tmp2485;
    wire tmp2486;
    wire tmp2487;
    wire tmp2488;
    wire tmp2489;
    wire tmp2490;
    wire tmp2491;
    wire tmp2492;
    wire tmp2493;
    wire tmp2494;
    wire tmp2495;
    wire tmp2496;
    wire tmp2497;
    wire tmp2498;
    wire tmp2499;
    wire tmp2500;
    wire tmp2501;
    wire tmp2502;
    wire tmp2503;
    wire tmp2504;
    wire tmp2505;
    wire tmp2506;
    wire tmp2507;
    wire tmp2508;
    wire tmp2509;
    wire tmp2510;
    wire tmp2511;
    wire tmp2512;
    wire tmp2513;
    wire tmp2514;
    wire tmp2515;
    wire tmp2516;
    wire tmp2517;
    wire tmp2518;
    wire tmp2519;
    wire tmp2520;
    wire tmp2521;
    wire tmp2522;
    wire tmp2523;
    wire tmp2524;
    wire tmp2525;
    wire tmp2526;
    wire tmp2527;
    wire tmp2528;
    wire tmp2529;
    wire tmp2530;
    wire tmp2531;
    wire tmp2532;
    wire tmp2533;
    wire tmp2534;
    wire tmp2535;
    wire tmp2536;
    wire tmp2537;
    wire tmp2538;
    wire tmp2539;
    wire tmp2540;
    wire tmp2541;
    wire tmp2542;
    wire tmp2543;
    wire tmp2544;
    wire tmp2545;
    wire tmp2546;
    wire tmp2547;
    wire tmp2548;
    wire tmp2549;
    wire tmp2550;
    wire tmp2551;
    wire tmp2552;
    wire tmp2553;
    wire tmp2554;
    wire tmp2555;
    wire tmp2556;
    wire tmp2557;
    wire tmp2558;
    wire tmp2559;
    wire tmp2560;
    wire tmp2561;
    wire tmp2562;
    wire tmp2563;
    wire tmp2564;
    wire tmp2565;
    wire tmp2566;
    wire tmp2567;
    wire tmp2568;
    wire[254:0] tmp2569;
    wire[255:0] tmp2570;
    wire tmp2571;
    wire[254:0] tmp2572;
    wire[255:0] tmp2573;
    wire tmp2574;
    wire tmp2575;
    wire[254:0] tmp2576;
    wire[255:0] tmp2577;
    wire tmp2578;
    wire tmp2579;
    wire[254:0] tmp2580;
    wire[255:0] tmp2581;
    wire tmp2582;
    wire tmp2583;
    wire tmp2584;
    wire tmp2585;
    wire tmp2586;
    wire tmp2587;
    wire tmp2588;
    wire tmp2589;
    wire tmp2590;
    wire tmp2591;
    wire tmp2592;
    wire tmp2593;
    wire tmp2594;
    wire tmp2595;
    wire tmp2596;
    wire tmp2597;
    wire tmp2598;
    wire tmp2599;
    wire tmp2600;
    wire tmp2601;
    wire tmp2602;
    wire tmp2603;
    wire[254:0] tmp2604;
    wire[255:0] tmp2605;
    wire[256:0] tmp2606;
    wire tmp2607;
    wire tmp2608;
    wire tmp2609;
    wire tmp2610;
    wire tmp2611;
    wire tmp2612;
    wire tmp2613;
    wire tmp2614;
    wire tmp2615;
    wire[254:0] tmp2616;
    wire[255:0] tmp2617;
    wire[256:0] tmp2618;
    wire tmp2619;
    wire tmp2620;
    wire tmp2621;
    wire tmp2622;
    wire tmp2623;
    wire tmp2624;
    wire tmp2625;
    wire tmp2626;
    wire tmp2627;
    wire tmp2628;
    wire tmp2629;
    wire tmp2630;
    wire tmp2631;
    wire tmp2632;
    wire tmp2633;
    wire tmp2634;
    wire tmp2635;
    wire tmp2636;
    wire tmp2637;
    wire tmp2638;
    wire tmp2639;
    wire tmp2640;
    wire tmp2641;
    wire tmp2642;
    wire tmp2643;
    wire tmp2644;
    wire tmp2645;
    wire tmp2646;
    wire tmp2647;
    wire tmp2648;
    wire tmp2649;
    wire tmp2650;
    wire tmp2651;
    wire tmp2652;
    wire[254:0] tmp2653;
    wire[255:0] tmp2654;
    wire[256:0] tmp2655;
    wire[1:0] tmp2656;
    wire[256:0] tmp2657;
    wire[256:0] tmp2658;
    wire[255:0] tmp2659;
    wire tmp2660;
    wire tmp2661;
    wire tmp2662;
    wire tmp2663;
    wire tmp2664;
    wire tmp2665;
    wire tmp2666;
    wire tmp2667;
    wire tmp2668;
    wire tmp2669;
    wire tmp2670;
    wire tmp2671;
    wire tmp2672;
    wire[254:0] tmp2673;
    wire[255:0] tmp2674;
    wire[256:0] tmp2675;
    wire[1:0] tmp2676;
    wire[256:0] tmp2677;
    wire[256:0] tmp2678;
    wire[255:0] tmp2679;
    wire tmp2680;
    wire tmp2681;
    wire tmp2682;
    wire tmp2683;
    wire tmp2684;
    wire tmp2685;
    wire tmp2686;
    wire tmp2687;
    wire tmp2688;
    wire tmp2689;
    wire tmp2690;
    wire tmp2691;
    wire tmp2692;
    wire[254:0] tmp2693;
    wire[255:0] tmp2694;
    wire[256:0] tmp2695;
    wire[1:0] tmp2696;
    wire[256:0] tmp2697;
    wire[256:0] tmp2698;
    wire[255:0] tmp2699;
    wire tmp2700;
    wire tmp2701;
    wire tmp2702;
    wire tmp2703;
    wire tmp2704;
    wire tmp2705;
    wire tmp2706;
    wire tmp2707;
    wire tmp2708;
    wire tmp2709;
    wire tmp2710;
    wire tmp2711;
    wire tmp2712;
    wire[254:0] tmp2713;
    wire[255:0] tmp2714;
    wire[256:0] tmp2715;
    wire[1:0] tmp2716;
    wire[256:0] tmp2717;
    wire[256:0] tmp2718;
    wire[255:0] tmp2719;
    wire tmp2720;
    wire tmp2721;
    wire tmp2722;
    wire tmp2723;
    wire tmp2724;
    wire tmp2725;
    wire tmp2726;
    wire tmp2727;
    wire tmp2728;
    wire tmp2729;
    wire tmp2730;
    wire tmp2731;
    wire[254:0] tmp2732;
    wire tmp2733;
    wire tmp2734;
    wire[255:0] tmp2735;
    wire tmp2736;
    wire tmp2737;
    wire[256:0] tmp2738;
    wire tmp2739;
    wire tmp2740;
    wire tmp2741;
    wire tmp2742;
    wire tmp2743;
    wire tmp2744;
    wire tmp2745;
    wire tmp2746;
    wire tmp2747;
    wire[254:0] tmp2748;
    wire tmp2749;
    wire tmp2750;
    wire[255:0] tmp2751;
    wire tmp2752;
    wire tmp2753;
    wire[256:0] tmp2754;
    wire tmp2755;
    wire tmp2756;
    wire tmp2757;
    wire tmp2758;
    wire tmp2759;
    wire tmp2760;
    wire tmp2761;
    wire tmp2762;
    wire tmp2763;
    wire tmp2764;
    wire[254:0] tmp2765;
    wire tmp2766;
    wire tmp2767;
    wire[255:0] tmp2768;
    wire tmp2769;
    wire tmp2770;
    wire[256:0] tmp2771;
    wire tmp2772;
    wire tmp2773;
    wire tmp2774;
    wire tmp2775;
    wire tmp2776;
    wire tmp2777;
    wire tmp2778;
    wire tmp2779;
    wire tmp2780;
    wire tmp2781;
    wire[254:0] tmp2782;
    wire tmp2783;
    wire tmp2784;
    wire[255:0] tmp2785;
    wire tmp2786;
    wire tmp2787;
    wire[256:0] tmp2788;
    wire tmp2789;
    wire tmp2790;
    wire tmp2791;
    wire tmp2792;
    wire tmp2793;
    wire tmp2794;
    wire tmp2795;
    wire tmp2796;
    wire tmp2797;
    wire tmp2798;
    wire tmp2799;
    wire tmp2800;
    wire tmp2801;
    wire tmp2802;
    wire tmp2803;
    wire tmp2804;
    wire tmp2805;
    wire tmp2806;
    wire tmp2807;
    wire tmp2808;
    wire tmp2809;
    wire tmp2810;
    wire tmp2811;
    wire tmp2812;
    wire tmp2813;
    wire tmp2814;
    wire tmp2815;
    wire tmp2816;
    wire tmp2817;
    wire tmp2818;
    wire tmp2819;
    wire tmp2820;
    wire tmp2821;
    wire tmp2822;
    wire tmp2823;
    wire tmp2824;
    wire tmp2825;
    wire tmp2826;
    wire[254:0] tmp2827;
    wire tmp2828;
    wire tmp2829;
    wire[255:0] tmp2830;
    wire tmp2831;
    wire tmp2832;
    wire tmp2833;
    wire tmp2834;
    wire tmp2835;
    wire tmp2836;
    wire tmp2837;
    wire tmp2838;
    wire tmp2839;
    wire tmp2840;
    wire tmp2841;
    wire tmp2842;
    wire tmp2843;
    wire tmp2844;
    wire tmp2845;
    wire[254:0] tmp2846;
    wire tmp2847;
    wire tmp2848;
    wire[255:0] tmp2849;
    wire tmp2850;
    wire tmp2851;
    wire tmp2852;
    wire tmp2853;
    wire tmp2854;
    wire tmp2855;
    wire tmp2856;
    wire tmp2857;
    wire tmp2858;
    wire tmp2859;
    wire tmp2860;
    wire tmp2861;
    wire tmp2862;
    wire tmp2863;
    wire tmp2864;
    wire[254:0] tmp2865;
    wire tmp2866;
    wire tmp2867;
    wire[255:0] tmp2868;
    wire tmp2869;
    wire tmp2870;
    wire tmp2871;
    wire tmp2872;
    wire tmp2873;
    wire tmp2874;
    wire tmp2875;
    wire tmp2876;
    wire tmp2877;
    wire tmp2878;
    wire tmp2879;
    wire tmp2880;
    wire tmp2881;
    wire tmp2882;
    wire tmp2883;
    wire[254:0] tmp2884;
    wire tmp2885;
    wire tmp2886;
    wire[255:0] tmp2887;
    wire tmp2888;
    wire tmp2889;
    wire tmp2890;
    wire tmp2891;
    wire tmp2892;
    wire tmp2893;
    wire tmp2894;
    wire tmp2895;
    wire tmp2896;
    wire tmp2897;
    wire tmp2898;
    wire tmp2899;
    wire tmp2900;
    wire tmp2901;
    wire tmp2902;
    wire tmp2903;
    wire tmp2904;
    wire tmp2905;
    wire tmp2906;
    wire tmp2907;
    wire tmp2908;
    wire tmp2909;
    wire tmp2910;
    wire tmp2911;
    wire tmp2912;
    wire tmp2913;
    wire tmp2914;
    wire tmp2915;
    wire tmp2916;
    wire tmp2917;
    wire tmp2918;
    wire tmp2919;
    wire tmp2920;
    wire tmp2921;
    wire tmp2922;
    wire tmp2923;
    wire tmp2924;
    wire tmp2925;
    wire tmp2926;
    wire tmp2927;
    wire tmp2928;
    wire tmp2929;
    wire tmp2930;
    wire tmp2931;
    wire tmp2932;
    wire tmp2933;
    wire tmp2934;
    wire tmp2935;
    wire tmp2936;
    wire tmp2937;
    wire tmp2938;
    wire tmp2939;
    wire tmp2940;
    wire tmp2941;
    wire tmp2942;
    wire tmp2943;
    wire tmp2944;
    wire tmp2945;
    wire tmp2946;
    wire tmp2947;
    wire tmp2948;
    wire tmp2949;
    wire tmp2950;
    wire tmp2951;
    wire tmp2952;
    wire tmp2953;
    wire tmp2954;
    wire tmp2955;
    wire tmp2956;
    wire tmp2957;
    wire tmp2958;
    wire tmp2959;
    wire tmp2960;
    wire tmp2961;
    wire tmp2962;
    wire tmp2963;
    wire tmp2964;
    wire tmp2965;
    wire tmp2966;
    wire tmp2967;
    wire tmp2968;
    wire tmp2969;
    wire tmp2970;
    wire tmp2971;
    wire tmp2972;
    wire tmp2973;
    wire tmp2974;
    wire tmp2975;
    wire tmp2976;
    wire tmp2977;
    wire tmp2978;
    wire tmp2979;
    wire tmp2980;
    wire tmp2981;
    wire tmp2982;
    wire tmp2983;
    wire tmp2984;
    wire tmp2985;
    wire tmp2986;
    wire tmp2987;
    wire tmp2988;
    wire tmp2989;
    wire tmp2990;
    wire tmp2991;
    wire tmp2992;
    wire tmp2993;
    wire tmp2994;
    wire tmp2995;
    wire tmp2996;
    wire tmp2997;
    wire tmp2998;
    wire tmp2999;
    wire tmp3000;
    wire tmp3001;
    wire tmp3002;
    wire tmp3003;
    wire tmp3004;
    wire tmp3005;
    wire tmp3006;
    wire tmp3007;
    wire tmp3008;
    wire tmp3009;
    wire tmp3010;
    wire tmp3011;
    wire tmp3012;
    wire tmp3013;
    wire tmp3014;
    wire tmp3015;
    wire tmp3016;
    wire tmp3017;
    wire tmp3018;
    wire tmp3019;
    wire tmp3020;
    wire tmp3021;
    wire tmp3022;
    wire tmp3023;
    wire tmp3024;
    wire tmp3025;
    wire tmp3026;
    wire[254:0] tmp3027;
    wire[255:0] tmp3028;
    wire tmp3029;
    wire[254:0] tmp3030;
    wire[255:0] tmp3031;
    wire tmp3032;
    wire[256:0] tmp3033;
    wire tmp3034;
    wire tmp3035;
    wire tmp3036;
    wire tmp3037;
    wire tmp3038;
    wire tmp3039;
    wire tmp3040;
    wire tmp3041;
    wire tmp3042;
    wire[254:0] tmp3043;
    wire[255:0] tmp3044;
    wire[256:0] tmp3045;
    wire tmp3046;
    wire tmp3047;
    wire tmp3048;
    wire tmp3049;
    wire tmp3050;
    wire tmp3051;
    wire tmp3052;
    wire tmp3053;
    wire tmp3054;
    wire tmp3055;
    wire[254:0] tmp3056;
    wire[255:0] tmp3057;
    wire[256:0] tmp3058;
    wire tmp3059;
    wire tmp3060;
    wire tmp3061;
    wire tmp3062;
    wire tmp3063;
    wire tmp3064;
    wire tmp3065;
    wire tmp3066;
    wire[254:0] tmp3067;
    wire[255:0] tmp3068;
    wire tmp3069;
    wire[256:0] tmp3070;
    wire tmp3071;
    wire tmp3072;
    wire tmp3073;
    wire tmp3074;
    wire tmp3075;
    wire tmp3076;
    wire tmp3077;
    wire tmp3078;
    wire tmp3079;
    wire tmp3080;
    wire[255:0] tmp3081;
    wire[255:0] tmp3082;
    wire tmp3083;
    wire tmp3084;
    wire tmp3085;
    wire tmp3086;
    wire tmp3087;
    wire tmp3088;
    wire tmp3089;
    wire tmp3090;
    wire tmp3091;
    wire tmp3092;
    wire tmp3093;
    wire tmp3094;
    wire tmp3095;
    wire tmp3096;
    wire tmp3097;
    wire tmp3098;
    wire[254:0] tmp3099;
    wire[255:0] tmp3100;
    wire tmp3101;
    wire[254:0] tmp3102;
    wire[255:0] tmp3103;
    wire tmp3104;
    wire[256:0] tmp3105;
    wire tmp3106;
    wire tmp3107;
    wire tmp3108;
    wire tmp3109;
    wire tmp3110;
    wire tmp3111;
    wire tmp3112;
    wire tmp3113;
    wire tmp3114;
    wire[254:0] tmp3115;
    wire[255:0] tmp3116;
    wire[256:0] tmp3117;
    wire tmp3118;
    wire tmp3119;
    wire tmp3120;
    wire tmp3121;
    wire tmp3122;
    wire tmp3123;
    wire tmp3124;
    wire tmp3125;
    wire tmp3126;
    wire tmp3127;
    wire[254:0] tmp3128;
    wire[255:0] tmp3129;
    wire[256:0] tmp3130;
    wire tmp3131;
    wire tmp3132;
    wire tmp3133;
    wire tmp3134;
    wire tmp3135;
    wire tmp3136;
    wire tmp3137;
    wire tmp3138;
    wire[254:0] tmp3139;
    wire[255:0] tmp3140;
    wire tmp3141;
    wire[256:0] tmp3142;
    wire tmp3143;
    wire tmp3144;
    wire tmp3145;
    wire tmp3146;
    wire tmp3147;
    wire tmp3148;
    wire tmp3149;
    wire tmp3150;
    wire tmp3151;
    wire tmp3152;
    wire[255:0] tmp3153;
    wire[255:0] tmp3154;
    wire tmp3155;
    wire tmp3156;
    wire tmp3157;
    wire tmp3158;
    wire tmp3159;
    wire tmp3160;
    wire tmp3161;
    wire tmp3162;
    wire tmp3163;
    wire tmp3164;
    wire tmp3165;
    wire tmp3166;
    wire tmp3167;
    wire tmp3168;
    wire tmp3169;
    wire tmp3170;
    wire[254:0] tmp3171;
    wire[255:0] tmp3172;
    wire tmp3173;
    wire[254:0] tmp3174;
    wire[255:0] tmp3175;
    wire tmp3176;
    wire[256:0] tmp3177;
    wire tmp3178;
    wire tmp3179;
    wire tmp3180;
    wire tmp3181;
    wire tmp3182;
    wire tmp3183;
    wire tmp3184;
    wire tmp3185;
    wire tmp3186;
    wire[254:0] tmp3187;
    wire[255:0] tmp3188;
    wire[256:0] tmp3189;
    wire tmp3190;
    wire tmp3191;
    wire tmp3192;
    wire tmp3193;
    wire tmp3194;
    wire tmp3195;
    wire tmp3196;
    wire tmp3197;
    wire tmp3198;
    wire tmp3199;
    wire[254:0] tmp3200;
    wire[255:0] tmp3201;
    wire[256:0] tmp3202;
    wire tmp3203;
    wire tmp3204;
    wire tmp3205;
    wire tmp3206;
    wire tmp3207;
    wire tmp3208;
    wire tmp3209;
    wire tmp3210;
    wire[254:0] tmp3211;
    wire[255:0] tmp3212;
    wire tmp3213;
    wire[256:0] tmp3214;
    wire tmp3215;
    wire tmp3216;
    wire tmp3217;
    wire tmp3218;
    wire tmp3219;
    wire tmp3220;
    wire tmp3221;
    wire tmp3222;
    wire tmp3223;
    wire tmp3224;
    wire[255:0] tmp3225;
    wire[255:0] tmp3226;
    wire tmp3227;
    wire tmp3228;
    wire tmp3229;
    wire tmp3230;
    wire tmp3231;
    wire tmp3232;
    wire tmp3233;
    wire tmp3234;
    wire tmp3235;
    wire tmp3236;
    wire tmp3237;
    wire tmp3238;
    wire tmp3239;
    wire tmp3240;
    wire tmp3241;
    wire tmp3242;
    wire[254:0] tmp3243;
    wire[255:0] tmp3244;
    wire tmp3245;
    wire[254:0] tmp3246;
    wire[255:0] tmp3247;
    wire tmp3248;
    wire[256:0] tmp3249;
    wire tmp3250;
    wire tmp3251;
    wire tmp3252;
    wire tmp3253;
    wire tmp3254;
    wire tmp3255;
    wire tmp3256;
    wire tmp3257;
    wire tmp3258;
    wire[254:0] tmp3259;
    wire[255:0] tmp3260;
    wire[256:0] tmp3261;
    wire tmp3262;
    wire tmp3263;
    wire tmp3264;
    wire tmp3265;
    wire tmp3266;
    wire tmp3267;
    wire tmp3268;
    wire tmp3269;
    wire tmp3270;
    wire tmp3271;
    wire[254:0] tmp3272;
    wire[255:0] tmp3273;
    wire[256:0] tmp3274;
    wire tmp3275;
    wire tmp3276;
    wire tmp3277;
    wire tmp3278;
    wire tmp3279;
    wire tmp3280;
    wire tmp3281;
    wire tmp3282;
    wire[254:0] tmp3283;
    wire[255:0] tmp3284;
    wire tmp3285;
    wire[256:0] tmp3286;
    wire tmp3287;
    wire tmp3288;
    wire tmp3289;
    wire tmp3290;
    wire tmp3291;
    wire tmp3292;
    wire tmp3293;
    wire tmp3294;
    wire tmp3295;
    wire tmp3296;
    wire[255:0] tmp3297;
    wire[255:0] tmp3298;
    wire tmp3299;
    wire tmp3300;
    wire tmp3301;
    wire tmp3302;
    wire tmp3303;
    wire tmp3304;
    wire tmp3305;
    wire tmp3306;
    wire tmp3307;
    wire tmp3308;
    wire tmp3309;
    wire tmp3310;
    wire tmp3311;
    wire tmp3312;
    wire tmp3313;
    wire tmp3314;
    wire tmp3315;
    wire tmp3316;
    wire[256:0] tmp3317;
    wire tmp3318;
    wire tmp3319;
    wire tmp3320;
    wire tmp3321;
    wire tmp3322;
    wire tmp3323;
    wire tmp3324;
    wire tmp3325;
    wire tmp3326;
    wire tmp3327;
    wire tmp3328;
    wire[256:0] tmp3329;
    wire tmp3330;
    wire tmp3331;
    wire tmp3332;
    wire tmp3333;
    wire tmp3334;
    wire tmp3335;
    wire tmp3336;
    wire tmp3337;
    wire tmp3338;
    wire tmp3339;
    wire tmp3340;
    wire tmp3341;
    wire[256:0] tmp3342;
    wire tmp3343;
    wire tmp3344;
    wire tmp3345;
    wire tmp3346;
    wire tmp3347;
    wire tmp3348;
    wire tmp3349;
    wire tmp3350;
    wire tmp3351;
    wire tmp3352;
    wire tmp3353;
    wire tmp3354;
    wire[256:0] tmp3355;
    wire tmp3356;
    wire tmp3357;
    wire tmp3358;
    wire tmp3359;
    wire tmp3360;
    wire tmp3361;
    wire tmp3362;
    wire tmp3363;
    wire tmp3364;
    wire tmp3365;
    wire[254:0] tmp3366;
    wire tmp3367;
    wire tmp3368;
    wire[255:0] tmp3369;
    wire tmp3370;
    wire tmp3371;
    wire[256:0] tmp3372;
    wire tmp3373;
    wire tmp3374;
    wire tmp3375;
    wire tmp3376;
    wire tmp3377;
    wire tmp3378;
    wire tmp3379;
    wire tmp3380;
    wire[254:0] tmp3381;
    wire tmp3382;
    wire tmp3383;
    wire[255:0] tmp3384;
    wire tmp3385;
    wire tmp3386;
    wire[256:0] tmp3387;
    wire tmp3388;
    wire tmp3389;
    wire tmp3390;
    wire tmp3391;
    wire tmp3392;
    wire tmp3393;
    wire tmp3394;
    wire tmp3395;
    wire[254:0] tmp3396;
    wire tmp3397;
    wire tmp3398;
    wire[255:0] tmp3399;
    wire tmp3400;
    wire tmp3401;
    wire[256:0] tmp3402;
    wire tmp3403;
    wire tmp3404;
    wire tmp3405;
    wire tmp3406;
    wire tmp3407;
    wire tmp3408;
    wire tmp3409;
    wire tmp3410;
    wire[254:0] tmp3411;
    wire tmp3412;
    wire tmp3413;
    wire[255:0] tmp3414;
    wire tmp3415;
    wire tmp3416;
    wire[256:0] tmp3417;
    wire tmp3418;
    wire tmp3419;
    wire tmp3420;
    wire tmp3421;
    wire tmp3422;
    wire tmp3423;
    wire tmp3424;
    wire tmp3425;
    wire tmp3426;
    wire tmp3427;
    wire tmp3428;
    wire tmp3429;
    wire tmp3430;
    wire tmp3431;
    wire tmp3432;
    wire tmp3433;
    wire tmp3434;
    wire tmp3435;
    wire tmp3436;
    wire tmp3437;
    wire tmp3438;
    wire tmp3439;
    wire tmp3440;
    wire tmp3441;
    wire tmp3442;
    wire tmp3443;
    wire tmp3444;
    wire tmp3445;
    wire tmp3446;
    wire tmp3447;
    wire tmp3448;
    wire tmp3449;
    wire tmp3450;
    wire tmp3451;
    wire tmp3452;
    wire tmp3453;
    wire tmp3454;
    wire tmp3455;
    wire tmp3456;
    wire tmp3457;
    wire tmp3458;
    wire tmp3459;
    wire tmp3460;
    wire tmp3461;
    wire tmp3462;
    wire tmp3463;
    wire tmp3464;
    wire tmp3465;
    wire tmp3466;
    wire tmp3467;
    wire tmp3468;
    wire tmp3469;
    wire tmp3470;
    wire tmp3471;
    wire tmp3472;
    wire tmp3473;
    wire tmp3474;
    wire[254:0] tmp3475;
    wire[255:0] tmp3476;
    wire[256:0] tmp3477;
    wire[1:0] tmp3478;
    wire[256:0] tmp3479;
    wire[256:0] tmp3480;
    wire tmp3481;
    wire[1:0] tmp3482;
    wire[257:0] tmp3483;
    wire tmp3484;
    wire tmp3485;
    wire[257:0] tmp3486;
    wire[258:0] tmp3487;
    wire[257:0] tmp3488;
    wire[255:0] tmp3489;
    wire tmp3490;
    wire[254:0] tmp3491;
    wire[255:0] tmp3492;
    wire tmp3493;
    wire[256:0] tmp3494;
    wire tmp3495;
    wire tmp3496;
    wire tmp3497;
    wire tmp3498;
    wire tmp3499;
    wire tmp3500;
    wire tmp3501;
    wire tmp3502;
    wire[255:0] tmp3503;
    wire[256:0] tmp3504;
    wire tmp3505;
    wire[257:0] tmp3506;
    wire tmp3507;
    wire tmp3508;
    wire tmp3509;
    wire tmp3510;
    wire tmp3511;
    wire tmp3512;
    wire tmp3513;
    wire tmp3514;
    wire tmp3515;
    wire tmp3516;
    wire[254:0] tmp3517;
    wire[255:0] tmp3518;
    wire[256:0] tmp3519;
    wire tmp3520;
    wire tmp3521;
    wire tmp3522;
    wire tmp3523;
    wire tmp3524;
    wire tmp3525;
    wire tmp3526;
    wire tmp3527;
    wire tmp3528;
    wire tmp3529;
    wire tmp3530;
    wire tmp3531;
    wire[254:0] tmp3532;
    wire[255:0] tmp3533;
    wire[256:0] tmp3534;
    wire tmp3535;
    wire tmp3536;
    wire tmp3537;
    wire tmp3538;
    wire tmp3539;
    wire tmp3540;
    wire tmp3541;
    wire tmp3542;
    wire tmp3543;
    wire[255:0] tmp3544;
    wire[256:0] tmp3545;
    wire[257:0] tmp3546;
    wire tmp3547;
    wire tmp3548;
    wire tmp3549;
    wire tmp3550;
    wire tmp3551;
    wire tmp3552;
    wire tmp3553;
    wire tmp3554;
    wire tmp3555;
    wire[254:0] tmp3556;
    wire[255:0] tmp3557;
    wire tmp3558;
    wire[256:0] tmp3559;
    wire tmp3560;
    wire tmp3561;
    wire tmp3562;
    wire tmp3563;
    wire tmp3564;
    wire tmp3565;
    wire tmp3566;
    wire tmp3567;
    wire tmp3568;
    wire tmp3569;
    wire[255:0] tmp3570;
    wire[255:0] tmp3571;
    wire tmp3572;
    wire tmp3573;
    wire tmp3574;
    wire tmp3575;
    wire tmp3576;
    wire tmp3577;
    wire tmp3578;
    wire tmp3579;
    wire tmp3580;
    wire tmp3581;
    wire tmp3582;
    wire tmp3583;
    wire tmp3584;
    wire tmp3585;
    wire tmp3586;
    wire tmp3587;
    wire tmp3588;
    wire tmp3589;
    wire tmp3590;
    wire tmp3591;
    wire tmp3592;
    wire tmp3593;
    wire tmp3594;
    wire tmp3595;
    wire tmp3596;
    wire tmp3597;
    wire tmp3598;
    wire tmp3599;
    wire tmp3600;
    wire tmp3601;
    wire tmp3602;
    wire tmp3603;
    wire tmp3604;
    wire[254:0] tmp3605;
    wire[255:0] tmp3606;
    wire[256:0] tmp3607;
    wire[1:0] tmp3608;
    wire[256:0] tmp3609;
    wire[256:0] tmp3610;
    wire tmp3611;
    wire[1:0] tmp3612;
    wire[257:0] tmp3613;
    wire tmp3614;
    wire tmp3615;
    wire[257:0] tmp3616;
    wire[258:0] tmp3617;
    wire[257:0] tmp3618;
    wire[255:0] tmp3619;
    wire tmp3620;
    wire[254:0] tmp3621;
    wire[255:0] tmp3622;
    wire tmp3623;
    wire[256:0] tmp3624;
    wire tmp3625;
    wire tmp3626;
    wire tmp3627;
    wire tmp3628;
    wire tmp3629;
    wire tmp3630;
    wire tmp3631;
    wire tmp3632;
    wire[255:0] tmp3633;
    wire[256:0] tmp3634;
    wire tmp3635;
    wire[257:0] tmp3636;
    wire tmp3637;
    wire tmp3638;
    wire tmp3639;
    wire tmp3640;
    wire tmp3641;
    wire tmp3642;
    wire tmp3643;
    wire tmp3644;
    wire tmp3645;
    wire tmp3646;
    wire[254:0] tmp3647;
    wire[255:0] tmp3648;
    wire[256:0] tmp3649;
    wire tmp3650;
    wire tmp3651;
    wire tmp3652;
    wire tmp3653;
    wire tmp3654;
    wire tmp3655;
    wire tmp3656;
    wire tmp3657;
    wire tmp3658;
    wire tmp3659;
    wire tmp3660;
    wire tmp3661;
    wire[254:0] tmp3662;
    wire[255:0] tmp3663;
    wire[256:0] tmp3664;
    wire tmp3665;
    wire tmp3666;
    wire tmp3667;
    wire tmp3668;
    wire tmp3669;
    wire tmp3670;
    wire tmp3671;
    wire tmp3672;
    wire tmp3673;
    wire[255:0] tmp3674;
    wire[256:0] tmp3675;
    wire[257:0] tmp3676;
    wire tmp3677;
    wire tmp3678;
    wire tmp3679;
    wire tmp3680;
    wire tmp3681;
    wire tmp3682;
    wire tmp3683;
    wire tmp3684;
    wire tmp3685;
    wire[254:0] tmp3686;
    wire[255:0] tmp3687;
    wire tmp3688;
    wire[256:0] tmp3689;
    wire tmp3690;
    wire tmp3691;
    wire tmp3692;
    wire tmp3693;
    wire tmp3694;
    wire tmp3695;
    wire tmp3696;
    wire tmp3697;
    wire tmp3698;
    wire tmp3699;
    wire[255:0] tmp3700;
    wire[255:0] tmp3701;
    wire tmp3702;
    wire tmp3703;
    wire tmp3704;
    wire tmp3705;
    wire tmp3706;
    wire tmp3707;
    wire tmp3708;
    wire tmp3709;
    wire tmp3710;
    wire tmp3711;
    wire tmp3712;
    wire tmp3713;
    wire tmp3714;
    wire tmp3715;
    wire tmp3716;
    wire tmp3717;
    wire tmp3718;
    wire tmp3719;
    wire tmp3720;
    wire tmp3721;
    wire tmp3722;
    wire tmp3723;
    wire tmp3724;
    wire tmp3725;
    wire tmp3726;
    wire tmp3727;
    wire tmp3728;
    wire tmp3729;
    wire tmp3730;
    wire tmp3731;
    wire tmp3732;
    wire tmp3733;
    wire tmp3734;
    wire[254:0] tmp3735;
    wire[255:0] tmp3736;
    wire[256:0] tmp3737;
    wire[1:0] tmp3738;
    wire[256:0] tmp3739;
    wire[256:0] tmp3740;
    wire tmp3741;
    wire[1:0] tmp3742;
    wire[257:0] tmp3743;
    wire tmp3744;
    wire tmp3745;
    wire[257:0] tmp3746;
    wire[258:0] tmp3747;
    wire[257:0] tmp3748;
    wire[255:0] tmp3749;
    wire tmp3750;
    wire[254:0] tmp3751;
    wire[255:0] tmp3752;
    wire tmp3753;
    wire[256:0] tmp3754;
    wire tmp3755;
    wire tmp3756;
    wire tmp3757;
    wire tmp3758;
    wire tmp3759;
    wire tmp3760;
    wire tmp3761;
    wire tmp3762;
    wire[255:0] tmp3763;
    wire[256:0] tmp3764;
    wire tmp3765;
    wire[257:0] tmp3766;
    wire tmp3767;
    wire tmp3768;
    wire tmp3769;
    wire tmp3770;
    wire tmp3771;
    wire tmp3772;
    wire tmp3773;
    wire tmp3774;
    wire tmp3775;
    wire tmp3776;
    wire[254:0] tmp3777;
    wire[255:0] tmp3778;
    wire[256:0] tmp3779;
    wire tmp3780;
    wire tmp3781;
    wire tmp3782;
    wire tmp3783;
    wire tmp3784;
    wire tmp3785;
    wire tmp3786;
    wire tmp3787;
    wire tmp3788;
    wire tmp3789;
    wire tmp3790;
    wire tmp3791;
    wire[254:0] tmp3792;
    wire[255:0] tmp3793;
    wire[256:0] tmp3794;
    wire tmp3795;
    wire tmp3796;
    wire tmp3797;
    wire tmp3798;
    wire tmp3799;
    wire tmp3800;
    wire tmp3801;
    wire tmp3802;
    wire tmp3803;
    wire[255:0] tmp3804;
    wire[256:0] tmp3805;
    wire[257:0] tmp3806;
    wire tmp3807;
    wire tmp3808;
    wire tmp3809;
    wire tmp3810;
    wire tmp3811;
    wire tmp3812;
    wire tmp3813;
    wire tmp3814;
    wire tmp3815;
    wire[254:0] tmp3816;
    wire[255:0] tmp3817;
    wire tmp3818;
    wire[256:0] tmp3819;
    wire tmp3820;
    wire tmp3821;
    wire tmp3822;
    wire tmp3823;
    wire tmp3824;
    wire tmp3825;
    wire tmp3826;
    wire tmp3827;
    wire tmp3828;
    wire tmp3829;
    wire[255:0] tmp3830;
    wire[255:0] tmp3831;
    wire tmp3832;
    wire tmp3833;
    wire tmp3834;
    wire tmp3835;
    wire tmp3836;
    wire tmp3837;
    wire tmp3838;
    wire tmp3839;
    wire tmp3840;
    wire tmp3841;
    wire tmp3842;
    wire tmp3843;
    wire tmp3844;
    wire tmp3845;
    wire tmp3846;
    wire tmp3847;
    wire tmp3848;
    wire tmp3849;
    wire tmp3850;
    wire tmp3851;
    wire tmp3852;
    wire tmp3853;
    wire tmp3854;
    wire tmp3855;
    wire tmp3856;
    wire tmp3857;
    wire tmp3858;
    wire tmp3859;
    wire tmp3860;
    wire tmp3861;
    wire tmp3862;
    wire tmp3863;
    wire tmp3864;
    wire[254:0] tmp3865;
    wire[255:0] tmp3866;
    wire[256:0] tmp3867;
    wire[1:0] tmp3868;
    wire[256:0] tmp3869;
    wire[256:0] tmp3870;
    wire tmp3871;
    wire[1:0] tmp3872;
    wire[257:0] tmp3873;
    wire tmp3874;
    wire tmp3875;
    wire[257:0] tmp3876;
    wire[258:0] tmp3877;
    wire[257:0] tmp3878;
    wire[255:0] tmp3879;
    wire tmp3880;
    wire[254:0] tmp3881;
    wire[255:0] tmp3882;
    wire tmp3883;
    wire[256:0] tmp3884;
    wire tmp3885;
    wire tmp3886;
    wire tmp3887;
    wire tmp3888;
    wire tmp3889;
    wire tmp3890;
    wire tmp3891;
    wire tmp3892;
    wire[255:0] tmp3893;
    wire[256:0] tmp3894;
    wire tmp3895;
    wire[257:0] tmp3896;
    wire tmp3897;
    wire tmp3898;
    wire tmp3899;
    wire tmp3900;
    wire tmp3901;
    wire tmp3902;
    wire tmp3903;
    wire tmp3904;
    wire tmp3905;
    wire tmp3906;
    wire[254:0] tmp3907;
    wire[255:0] tmp3908;
    wire[256:0] tmp3909;
    wire tmp3910;
    wire tmp3911;
    wire tmp3912;
    wire tmp3913;
    wire tmp3914;
    wire tmp3915;
    wire tmp3916;
    wire tmp3917;
    wire tmp3918;
    wire tmp3919;
    wire tmp3920;
    wire tmp3921;
    wire[254:0] tmp3922;
    wire[255:0] tmp3923;
    wire[256:0] tmp3924;
    wire tmp3925;
    wire tmp3926;
    wire tmp3927;
    wire tmp3928;
    wire tmp3929;
    wire tmp3930;
    wire tmp3931;
    wire tmp3932;
    wire tmp3933;
    wire[255:0] tmp3934;
    wire[256:0] tmp3935;
    wire[257:0] tmp3936;
    wire tmp3937;
    wire tmp3938;
    wire tmp3939;
    wire tmp3940;
    wire tmp3941;
    wire tmp3942;
    wire tmp3943;
    wire tmp3944;
    wire tmp3945;
    wire[254:0] tmp3946;
    wire[255:0] tmp3947;
    wire tmp3948;
    wire[256:0] tmp3949;
    wire tmp3950;
    wire tmp3951;
    wire tmp3952;
    wire tmp3953;
    wire tmp3954;
    wire tmp3955;
    wire tmp3956;
    wire tmp3957;
    wire tmp3958;
    wire tmp3959;
    wire[255:0] tmp3960;
    wire[255:0] tmp3961;
    wire tmp3962;
    wire tmp3963;
    wire tmp3964;
    wire tmp3965;
    wire tmp3966;
    wire tmp3967;
    wire tmp3968;
    wire tmp3969;
    wire tmp3970;
    wire tmp3971;
    wire tmp3972;
    wire tmp3973;
    wire tmp3974;
    wire tmp3975;
    wire tmp3976;
    wire tmp3977;
    wire tmp3978;
    wire tmp3979;
    wire[256:0] tmp3980;
    wire tmp3981;
    wire tmp3982;
    wire tmp3983;
    wire tmp3984;
    wire tmp3985;
    wire tmp3986;
    wire tmp3987;
    wire tmp3988;
    wire tmp3989;
    wire[256:0] tmp3990;
    wire tmp3991;
    wire tmp3992;
    wire tmp3993;
    wire tmp3994;
    wire tmp3995;
    wire tmp3996;
    wire tmp3997;
    wire tmp3998;
    wire tmp3999;
    wire tmp4000;
    wire[256:0] tmp4001;
    wire tmp4002;
    wire tmp4003;
    wire tmp4004;
    wire tmp4005;
    wire tmp4006;
    wire tmp4007;
    wire tmp4008;
    wire tmp4009;
    wire tmp4010;
    wire tmp4011;
    wire[256:0] tmp4012;
    wire tmp4013;
    wire tmp4014;
    wire tmp4015;
    wire tmp4016;
    wire tmp4017;
    wire tmp4018;
    wire tmp4019;
    wire tmp4020;
    wire tmp4021;
    wire tmp4022;
    wire tmp4023;
    wire tmp4024;
    wire tmp4025;
    wire tmp4026;
    wire tmp4027;
    wire tmp4028;
    wire tmp4029;
    wire tmp4030;
    wire tmp4031;
    wire tmp4032;
    wire tmp4033;
    wire tmp4034;
    wire tmp4035;
    wire tmp4036;
    wire tmp4037;
    wire tmp4038;
    wire tmp4039;
    wire tmp4040;
    wire tmp4041;
    wire tmp4042;
    wire tmp4043;
    wire tmp4044;
    wire tmp4045;
    wire tmp4046;
    wire tmp4047;
    wire tmp4048;
    wire tmp4049;
    wire tmp4050;
    wire tmp4051;
    wire tmp4052;
    wire tmp4053;
    wire tmp4054;
    wire tmp4055;
    wire tmp4056;
    wire tmp4057;
    wire tmp4058;
    wire tmp4059;
    wire tmp4060;
    wire tmp4061;
    wire tmp4062;
    wire tmp4063;
    wire tmp4064;
    wire tmp4065;
    wire tmp4066;
    wire tmp4067;
    wire tmp4068;
    wire tmp4069;
    wire tmp4070;
    wire tmp4071;
    wire tmp4072;
    wire tmp4073;
    wire tmp4074;
    wire tmp4075;
    wire tmp4076;
    wire tmp4077;
    wire tmp4078;
    wire tmp4079;
    wire tmp4080;
    wire tmp4081;
    wire tmp4082;
    wire tmp4083;
    wire tmp4084;
    wire tmp4085;
    wire tmp4086;
    wire tmp4087;
    wire tmp4088;
    wire tmp4089;
    wire tmp4090;
    wire tmp4091;
    wire tmp4092;
    wire tmp4093;
    wire tmp4094;
    wire tmp4095;
    wire tmp4096;
    wire tmp4097;
    wire tmp4098;
    wire tmp4099;
    wire tmp4100;
    wire tmp4101;
    wire tmp4102;
    wire tmp4103;
    wire tmp4104;
    wire tmp4105;
    wire tmp4106;
    wire tmp4107;
    wire tmp4108;
    wire tmp4109;
    wire tmp4110;
    wire tmp4111;
    wire tmp4112;
    wire tmp4113;
    wire tmp4114;
    wire tmp4115;
    wire tmp4116;
    wire tmp4117;
    wire tmp4118;
    wire tmp4119;
    wire tmp4120;
    wire tmp4121;
    wire tmp4122;
    wire tmp4123;
    wire tmp4124;
    wire tmp4125;
    wire tmp4126;
    wire tmp4127;
    wire tmp4128;
    wire tmp4129;
    wire tmp4130;
    wire tmp4131;
    wire tmp4132;
    wire tmp4133;
    wire tmp4134;
    wire tmp4135;
    wire tmp4136;
    wire tmp4137;
    wire tmp4138;
    wire tmp4139;
    wire tmp4140;
    wire tmp4141;
    wire tmp4142;
    wire tmp4143;
    wire tmp4144;
    wire tmp4145;
    wire tmp4146;
    wire tmp4147;
    wire tmp4148;
    wire tmp4149;
    wire tmp4150;
    wire tmp4151;
    wire tmp4152;
    wire tmp4153;
    wire tmp4154;
    wire tmp4155;
    wire tmp4156;
    wire tmp4157;
    wire tmp4158;
    wire tmp4159;
    wire tmp4160;
    wire tmp4161;
    wire tmp4162;
    wire tmp4163;
    wire tmp4164;
    wire tmp4165;
    wire tmp4166;
    wire tmp4167;
    wire tmp4168;
    wire tmp4169;
    wire tmp4170;
    wire tmp4171;
    wire tmp4172;
    wire tmp4173;
    wire tmp4174;
    wire tmp4175;
    wire tmp4176;
    wire tmp4177;
    wire tmp4178;
    wire tmp4179;
    wire tmp4180;
    wire tmp4181;
    wire tmp4182;
    wire tmp4183;
    wire tmp4184;
    wire tmp4185;
    wire tmp4186;
    wire tmp4187;
    wire tmp4188;
    wire tmp4189;
    wire tmp4190;
    wire tmp4191;
    wire tmp4192;
    wire tmp4193;
    wire tmp4194;
    wire tmp4195;
    wire tmp4196;
    wire tmp4197;
    wire tmp4198;
    wire tmp4199;
    wire tmp4200;
    wire tmp4201;
    wire tmp4202;
    wire[256:0] tmp4203;
    wire tmp4204;
    wire tmp4205;
    wire tmp4206;
    wire tmp4207;
    wire tmp4208;
    wire tmp4209;
    wire tmp4210;
    wire[253:0] tmp4211;
    wire[255:0] tmp4212;
    wire tmp4213;
    wire[254:0] tmp4214;
    wire[255:0] tmp4215;
    wire tmp4216;
    wire[256:0] tmp4217;
    wire tmp4218;
    wire tmp4219;
    wire tmp4220;
    wire tmp4221;
    wire tmp4222;
    wire tmp4223;
    wire tmp4224;
    wire tmp4225;
    wire tmp4226;
    wire[254:0] tmp4227;
    wire[255:0] tmp4228;
    wire[256:0] tmp4229;
    wire tmp4230;
    wire tmp4231;
    wire tmp4232;
    wire tmp4233;
    wire tmp4234;
    wire tmp4235;
    wire tmp4236;
    wire tmp4237;
    wire tmp4238;
    wire tmp4239;
    wire[254:0] tmp4240;
    wire[255:0] tmp4241;
    wire[256:0] tmp4242;
    wire tmp4243;
    wire tmp4244;
    wire tmp4245;
    wire tmp4246;
    wire tmp4247;
    wire tmp4248;
    wire tmp4249;
    wire tmp4250;
    wire[254:0] tmp4251;
    wire[255:0] tmp4252;
    wire tmp4253;
    wire[256:0] tmp4254;
    wire tmp4255;
    wire tmp4256;
    wire tmp4257;
    wire tmp4258;
    wire tmp4259;
    wire tmp4260;
    wire tmp4261;
    wire tmp4262;
    wire tmp4263;
    wire tmp4264;
    wire[255:0] tmp4265;
    wire[255:0] tmp4266;
    wire tmp4267;
    wire tmp4268;
    wire[256:0] tmp4269;
    wire tmp4270;
    wire tmp4271;
    wire tmp4272;
    wire tmp4273;
    wire tmp4274;
    wire tmp4275;
    wire tmp4276;
    wire tmp4277;
    wire tmp4278;
    wire tmp4279;
    wire[256:0] tmp4280;
    wire tmp4281;
    wire tmp4282;
    wire tmp4283;
    wire tmp4284;
    wire tmp4285;
    wire tmp4286;
    wire tmp4287;
    wire tmp4288;
    wire[253:0] tmp4289;
    wire[255:0] tmp4290;
    wire tmp4291;
    wire[254:0] tmp4292;
    wire[255:0] tmp4293;
    wire tmp4294;
    wire[256:0] tmp4295;
    wire tmp4296;
    wire tmp4297;
    wire tmp4298;
    wire tmp4299;
    wire tmp4300;
    wire tmp4301;
    wire tmp4302;
    wire tmp4303;
    wire tmp4304;
    wire[254:0] tmp4305;
    wire[255:0] tmp4306;
    wire[256:0] tmp4307;
    wire tmp4308;
    wire tmp4309;
    wire tmp4310;
    wire tmp4311;
    wire tmp4312;
    wire tmp4313;
    wire tmp4314;
    wire tmp4315;
    wire tmp4316;
    wire tmp4317;
    wire[254:0] tmp4318;
    wire[255:0] tmp4319;
    wire[256:0] tmp4320;
    wire tmp4321;
    wire tmp4322;
    wire tmp4323;
    wire tmp4324;
    wire tmp4325;
    wire tmp4326;
    wire tmp4327;
    wire tmp4328;
    wire[254:0] tmp4329;
    wire[255:0] tmp4330;
    wire tmp4331;
    wire[256:0] tmp4332;
    wire tmp4333;
    wire tmp4334;
    wire tmp4335;
    wire tmp4336;
    wire tmp4337;
    wire tmp4338;
    wire tmp4339;
    wire tmp4340;
    wire tmp4341;
    wire tmp4342;
    wire[255:0] tmp4343;
    wire[255:0] tmp4344;
    wire tmp4345;
    wire tmp4346;
    wire[256:0] tmp4347;
    wire tmp4348;
    wire tmp4349;
    wire tmp4350;
    wire tmp4351;
    wire tmp4352;
    wire tmp4353;
    wire tmp4354;
    wire tmp4355;
    wire tmp4356;
    wire tmp4357;
    wire[256:0] tmp4358;
    wire tmp4359;
    wire tmp4360;
    wire tmp4361;
    wire tmp4362;
    wire tmp4363;
    wire tmp4364;
    wire tmp4365;
    wire tmp4366;
    wire[253:0] tmp4367;
    wire[255:0] tmp4368;
    wire tmp4369;
    wire[254:0] tmp4370;
    wire[255:0] tmp4371;
    wire tmp4372;
    wire[256:0] tmp4373;
    wire tmp4374;
    wire tmp4375;
    wire tmp4376;
    wire tmp4377;
    wire tmp4378;
    wire tmp4379;
    wire tmp4380;
    wire tmp4381;
    wire tmp4382;
    wire[254:0] tmp4383;
    wire[255:0] tmp4384;
    wire[256:0] tmp4385;
    wire tmp4386;
    wire tmp4387;
    wire tmp4388;
    wire tmp4389;
    wire tmp4390;
    wire tmp4391;
    wire tmp4392;
    wire tmp4393;
    wire tmp4394;
    wire tmp4395;
    wire[254:0] tmp4396;
    wire[255:0] tmp4397;
    wire[256:0] tmp4398;
    wire tmp4399;
    wire tmp4400;
    wire tmp4401;
    wire tmp4402;
    wire tmp4403;
    wire tmp4404;
    wire tmp4405;
    wire tmp4406;
    wire[254:0] tmp4407;
    wire[255:0] tmp4408;
    wire tmp4409;
    wire[256:0] tmp4410;
    wire tmp4411;
    wire tmp4412;
    wire tmp4413;
    wire tmp4414;
    wire tmp4415;
    wire tmp4416;
    wire tmp4417;
    wire tmp4418;
    wire tmp4419;
    wire tmp4420;
    wire[255:0] tmp4421;
    wire[255:0] tmp4422;
    wire tmp4423;
    wire tmp4424;
    wire[256:0] tmp4425;
    wire tmp4426;
    wire tmp4427;
    wire tmp4428;
    wire tmp4429;
    wire tmp4430;
    wire tmp4431;
    wire tmp4432;
    wire tmp4433;
    wire tmp4434;
    wire tmp4435;
    wire[256:0] tmp4436;
    wire tmp4437;
    wire tmp4438;
    wire tmp4439;
    wire tmp4440;
    wire tmp4441;
    wire tmp4442;
    wire tmp4443;
    wire tmp4444;
    wire[253:0] tmp4445;
    wire[255:0] tmp4446;
    wire tmp4447;
    wire[254:0] tmp4448;
    wire[255:0] tmp4449;
    wire tmp4450;
    wire[256:0] tmp4451;
    wire tmp4452;
    wire tmp4453;
    wire tmp4454;
    wire tmp4455;
    wire tmp4456;
    wire tmp4457;
    wire tmp4458;
    wire tmp4459;
    wire tmp4460;
    wire[254:0] tmp4461;
    wire[255:0] tmp4462;
    wire[256:0] tmp4463;
    wire tmp4464;
    wire tmp4465;
    wire tmp4466;
    wire tmp4467;
    wire tmp4468;
    wire tmp4469;
    wire tmp4470;
    wire tmp4471;
    wire tmp4472;
    wire tmp4473;
    wire[254:0] tmp4474;
    wire[255:0] tmp4475;
    wire[256:0] tmp4476;
    wire tmp4477;
    wire tmp4478;
    wire tmp4479;
    wire tmp4480;
    wire tmp4481;
    wire tmp4482;
    wire tmp4483;
    wire tmp4484;
    wire[254:0] tmp4485;
    wire[255:0] tmp4486;
    wire tmp4487;
    wire[256:0] tmp4488;
    wire tmp4489;
    wire tmp4490;
    wire tmp4491;
    wire tmp4492;
    wire tmp4493;
    wire tmp4494;
    wire tmp4495;
    wire tmp4496;
    wire tmp4497;
    wire tmp4498;
    wire[255:0] tmp4499;
    wire[255:0] tmp4500;
    wire tmp4501;
    wire tmp4502;
    wire[256:0] tmp4503;
    wire tmp4504;
    wire tmp4505;
    wire tmp4506;
    wire tmp4507;
    wire tmp4508;
    wire tmp4509;
    wire tmp4510;
    wire tmp4511;
    wire tmp4512;
    wire tmp4513;
    wire tmp4514;
    wire tmp4515;
    wire tmp4516;
    wire tmp4517;
    wire tmp4518;
    wire tmp4519;
    wire tmp4520;
    wire tmp4521;
    wire tmp4522;
    wire tmp4523;
    wire tmp4524;
    wire tmp4525;
    wire tmp4526;
    wire tmp4527;
    wire tmp4528;
    wire tmp4529;
    wire tmp4530;
    wire tmp4531;
    wire tmp4532;
    wire tmp4533;
    wire tmp4534;
    wire tmp4535;
    wire tmp4536;
    wire tmp4537;
    wire tmp4538;
    wire tmp4539;
    wire tmp4540;
    wire tmp4541;
    wire tmp4542;
    wire tmp4543;
    wire tmp4544;
    wire tmp4545;
    wire tmp4546;
    wire tmp4547;
    wire tmp4548;
    wire tmp4549;
    wire tmp4550;
    wire tmp4551;
    wire tmp4552;
    wire tmp4553;
    wire[254:0] tmp4554;
    wire tmp4555;
    wire tmp4556;
    wire[255:0] tmp4557;
    wire tmp4558;
    wire tmp4559;
    wire tmp4560;
    wire tmp4561;
    wire tmp4562;
    wire tmp4563;
    wire tmp4564;
    wire tmp4565;
    wire tmp4566;
    wire tmp4567;
    wire tmp4568;
    wire tmp4569;
    wire tmp4570;
    wire tmp4571;
    wire tmp4572;
    wire tmp4573;
    wire tmp4574;
    wire tmp4575;
    wire tmp4576;
    wire tmp4577;
    wire tmp4578;
    wire tmp4579;
    wire[254:0] tmp4580;
    wire tmp4581;
    wire tmp4582;
    wire[255:0] tmp4583;
    wire tmp4584;
    wire tmp4585;
    wire tmp4586;
    wire tmp4587;
    wire tmp4588;
    wire tmp4589;
    wire tmp4590;
    wire tmp4591;
    wire tmp4592;
    wire tmp4593;
    wire tmp4594;
    wire tmp4595;
    wire tmp4596;
    wire tmp4597;
    wire tmp4598;
    wire tmp4599;
    wire tmp4600;
    wire tmp4601;
    wire tmp4602;
    wire tmp4603;
    wire tmp4604;
    wire tmp4605;
    wire[254:0] tmp4606;
    wire tmp4607;
    wire tmp4608;
    wire[255:0] tmp4609;
    wire tmp4610;
    wire tmp4611;
    wire tmp4612;
    wire tmp4613;
    wire tmp4614;
    wire tmp4615;
    wire tmp4616;
    wire tmp4617;
    wire tmp4618;
    wire tmp4619;
    wire tmp4620;
    wire tmp4621;
    wire tmp4622;
    wire tmp4623;
    wire tmp4624;
    wire tmp4625;
    wire tmp4626;
    wire tmp4627;
    wire tmp4628;
    wire tmp4629;
    wire tmp4630;
    wire tmp4631;
    wire[254:0] tmp4632;
    wire tmp4633;
    wire tmp4634;
    wire[255:0] tmp4635;
    wire tmp4636;
    wire tmp4637;
    wire tmp4638;
    wire tmp4639;
    wire tmp4640;
    wire tmp4641;
    wire tmp4642;
    wire tmp4643;
    wire tmp4644;
    wire tmp4645;
    wire tmp4646;
    wire tmp4647;
    wire tmp4648;
    wire tmp4649;
    wire tmp4650;
    wire tmp4651;
    wire tmp4652;
    wire tmp4653;
    wire tmp4654;
    wire tmp4655;
    wire tmp4656;
    wire tmp4657;
    wire tmp4658;
    wire tmp4659;
    wire tmp4660;
    wire tmp4661;
    wire tmp4662;
    wire tmp4663;
    wire tmp4664;
    wire tmp4665;
    wire tmp4666;
    wire tmp4667;
    wire tmp4668;
    wire tmp4669;
    wire tmp4670;
    wire tmp4671;
    wire tmp4672;
    wire tmp4673;
    wire tmp4674;
    wire tmp4675;
    wire tmp4676;
    wire tmp4677;
    wire tmp4678;
    wire tmp4679;
    wire tmp4680;
    wire tmp4681;
    wire tmp4682;
    wire tmp4683;
    wire tmp4684;
    wire tmp4685;
    wire tmp4686;
    wire tmp4687;
    wire tmp4688;
    wire tmp4689;
    wire tmp4690;
    wire tmp4691;
    wire tmp4692;
    wire tmp4693;
    wire tmp4694;
    wire tmp4695;
    wire tmp4696;
    wire tmp4697;
    wire tmp4698;
    wire tmp4699;
    wire tmp4700;
    wire tmp4701;
    wire tmp4702;
    wire tmp4703;
    wire tmp4704;
    wire tmp4705;
    wire tmp4706;
    wire tmp4707;
    wire tmp4708;
    wire tmp4709;
    wire tmp4710;
    wire tmp4711;
    wire tmp4712;
    wire tmp4713;
    wire tmp4714;
    wire tmp4715;
    wire tmp4716;
    wire tmp4717;
    wire tmp4718;
    wire tmp4719;
    wire tmp4720;
    wire tmp4721;
    wire tmp4722;
    wire tmp4723;
    wire tmp4724;
    wire tmp4725;
    wire tmp4726;
    wire tmp4727;
    wire tmp4728;
    wire tmp4729;
    wire tmp4730;
    wire tmp4731;
    wire tmp4732;
    wire tmp4733;
    wire tmp4734;
    wire tmp4735;
    wire tmp4736;
    wire tmp4737;
    wire tmp4738;
    wire tmp4739;
    wire tmp4740;
    wire tmp4741;
    wire tmp4742;
    wire tmp4743;
    wire tmp4744;
    wire tmp4745;
    wire tmp4746;
    wire tmp4747;
    wire tmp4748;
    wire tmp4749;
    wire tmp4750;
    wire tmp4751;
    wire tmp4752;
    wire tmp4753;
    wire tmp4754;
    wire tmp4755;
    wire tmp4756;
    wire tmp4757;
    wire tmp4758;
    wire tmp4759;
    wire tmp4760;
    wire tmp4761;
    wire tmp4762;
    wire tmp4763;
    wire tmp4764;
    wire tmp4765;
    wire tmp4766;
    wire tmp4767;
    wire tmp4768;
    wire tmp4769;
    wire tmp4770;
    wire tmp4771;
    wire tmp4772;
    wire tmp4773;
    wire tmp4774;
    wire tmp4775;
    wire tmp4776;
    wire tmp4777;
    wire tmp4778;
    wire tmp4779;
    wire tmp4780;
    wire tmp4781;
    wire tmp4782;
    wire tmp4783;
    wire tmp4784;
    wire tmp4785;
    wire tmp4786;
    wire tmp4787;
    wire tmp4788;
    wire tmp4789;
    wire tmp4790;
    wire tmp4791;
    wire tmp4792;
    wire tmp4793;
    wire tmp4794;
    wire tmp4795;
    wire tmp4796;
    wire tmp4797;
    wire tmp4798;
    wire tmp4799;
    wire tmp4800;
    wire tmp4801;
    wire tmp4802;
    wire tmp4803;
    wire tmp4804;
    wire tmp4805;
    wire tmp4806;
    wire tmp4807;
    wire tmp4808;
    wire tmp4809;
    wire tmp4810;
    wire tmp4811;
    wire tmp4812;
    wire tmp4813;
    wire tmp4814;
    wire tmp4815;
    wire tmp4816;
    wire tmp4817;
    wire tmp4818;
    wire tmp4819;
    wire tmp4820;
    wire tmp4821;
    wire tmp4822;
    wire tmp4823;
    wire tmp4824;
    wire tmp4825;
    wire tmp4826;
    wire tmp4827;
    wire tmp4828;
    wire tmp4829;
    wire tmp4830;
    wire tmp4831;
    wire tmp4832;
    wire tmp4833;
    wire tmp4834;
    wire tmp4835;
    wire tmp4836;
    wire tmp4837;
    wire[254:0] tmp4838;
    wire[255:0] tmp4839;
    wire tmp4840;
    wire[254:0] tmp4841;
    wire[255:0] tmp4842;
    wire tmp4843;
    wire[256:0] tmp4844;
    wire tmp4845;
    wire tmp4846;
    wire tmp4847;
    wire tmp4848;
    wire tmp4849;
    wire tmp4850;
    wire tmp4851;
    wire tmp4852;
    wire tmp4853;
    wire[254:0] tmp4854;
    wire[255:0] tmp4855;
    wire[256:0] tmp4856;
    wire tmp4857;
    wire tmp4858;
    wire tmp4859;
    wire tmp4860;
    wire tmp4861;
    wire tmp4862;
    wire tmp4863;
    wire tmp4864;
    wire tmp4865;
    wire tmp4866;
    wire[254:0] tmp4867;
    wire[255:0] tmp4868;
    wire[256:0] tmp4869;
    wire tmp4870;
    wire tmp4871;
    wire tmp4872;
    wire tmp4873;
    wire tmp4874;
    wire tmp4875;
    wire tmp4876;
    wire tmp4877;
    wire[254:0] tmp4878;
    wire[255:0] tmp4879;
    wire tmp4880;
    wire[256:0] tmp4881;
    wire tmp4882;
    wire tmp4883;
    wire tmp4884;
    wire tmp4885;
    wire tmp4886;
    wire tmp4887;
    wire tmp4888;
    wire tmp4889;
    wire tmp4890;
    wire tmp4891;
    wire[255:0] tmp4892;
    wire[255:0] tmp4893;
    wire tmp4894;
    wire tmp4895;
    wire tmp4896;
    wire tmp4897;
    wire tmp4898;
    wire tmp4899;
    wire tmp4900;
    wire tmp4901;
    wire tmp4902;
    wire tmp4903;
    wire tmp4904;
    wire tmp4905;
    wire tmp4906;
    wire tmp4907;
    wire tmp4908;
    wire tmp4909;
    wire tmp4910;
    wire tmp4911;
    wire tmp4912;
    wire tmp4913;
    wire tmp4914;
    wire tmp4915;
    wire tmp4916;
    wire[254:0] tmp4917;
    wire[255:0] tmp4918;
    wire tmp4919;
    wire[254:0] tmp4920;
    wire[255:0] tmp4921;
    wire tmp4922;
    wire[256:0] tmp4923;
    wire tmp4924;
    wire tmp4925;
    wire tmp4926;
    wire tmp4927;
    wire tmp4928;
    wire tmp4929;
    wire tmp4930;
    wire tmp4931;
    wire tmp4932;
    wire[254:0] tmp4933;
    wire[255:0] tmp4934;
    wire[256:0] tmp4935;
    wire tmp4936;
    wire tmp4937;
    wire tmp4938;
    wire tmp4939;
    wire tmp4940;
    wire tmp4941;
    wire tmp4942;
    wire tmp4943;
    wire tmp4944;
    wire tmp4945;
    wire[254:0] tmp4946;
    wire[255:0] tmp4947;
    wire[256:0] tmp4948;
    wire tmp4949;
    wire tmp4950;
    wire tmp4951;
    wire tmp4952;
    wire tmp4953;
    wire tmp4954;
    wire tmp4955;
    wire tmp4956;
    wire[254:0] tmp4957;
    wire[255:0] tmp4958;
    wire tmp4959;
    wire[256:0] tmp4960;
    wire tmp4961;
    wire tmp4962;
    wire tmp4963;
    wire tmp4964;
    wire tmp4965;
    wire tmp4966;
    wire tmp4967;
    wire tmp4968;
    wire tmp4969;
    wire tmp4970;
    wire[255:0] tmp4971;
    wire[255:0] tmp4972;
    wire tmp4973;
    wire tmp4974;
    wire tmp4975;
    wire tmp4976;
    wire tmp4977;
    wire tmp4978;
    wire tmp4979;
    wire tmp4980;
    wire tmp4981;
    wire tmp4982;
    wire tmp4983;
    wire tmp4984;
    wire tmp4985;
    wire tmp4986;
    wire tmp4987;
    wire tmp4988;
    wire tmp4989;
    wire tmp4990;
    wire tmp4991;
    wire tmp4992;
    wire tmp4993;
    wire tmp4994;
    wire tmp4995;
    wire[254:0] tmp4996;
    wire[255:0] tmp4997;
    wire tmp4998;
    wire[254:0] tmp4999;
    wire[255:0] tmp5000;
    wire tmp5001;
    wire[256:0] tmp5002;
    wire tmp5003;
    wire tmp5004;
    wire tmp5005;
    wire tmp5006;
    wire tmp5007;
    wire tmp5008;
    wire tmp5009;
    wire tmp5010;
    wire tmp5011;
    wire[254:0] tmp5012;
    wire[255:0] tmp5013;
    wire[256:0] tmp5014;
    wire tmp5015;
    wire tmp5016;
    wire tmp5017;
    wire tmp5018;
    wire tmp5019;
    wire tmp5020;
    wire tmp5021;
    wire tmp5022;
    wire tmp5023;
    wire tmp5024;
    wire[254:0] tmp5025;
    wire[255:0] tmp5026;
    wire[256:0] tmp5027;
    wire tmp5028;
    wire tmp5029;
    wire tmp5030;
    wire tmp5031;
    wire tmp5032;
    wire tmp5033;
    wire tmp5034;
    wire tmp5035;
    wire[254:0] tmp5036;
    wire[255:0] tmp5037;
    wire tmp5038;
    wire[256:0] tmp5039;
    wire tmp5040;
    wire tmp5041;
    wire tmp5042;
    wire tmp5043;
    wire tmp5044;
    wire tmp5045;
    wire tmp5046;
    wire tmp5047;
    wire tmp5048;
    wire tmp5049;
    wire[255:0] tmp5050;
    wire[255:0] tmp5051;
    wire tmp5052;
    wire tmp5053;
    wire tmp5054;
    wire tmp5055;
    wire tmp5056;
    wire tmp5057;
    wire tmp5058;
    wire tmp5059;
    wire tmp5060;
    wire tmp5061;
    wire tmp5062;
    wire tmp5063;
    wire tmp5064;
    wire tmp5065;
    wire tmp5066;
    wire tmp5067;
    wire tmp5068;
    wire tmp5069;
    wire tmp5070;
    wire tmp5071;
    wire tmp5072;
    wire tmp5073;
    wire tmp5074;
    wire[254:0] tmp5075;
    wire[255:0] tmp5076;
    wire tmp5077;
    wire[254:0] tmp5078;
    wire[255:0] tmp5079;
    wire tmp5080;
    wire[256:0] tmp5081;
    wire tmp5082;
    wire tmp5083;
    wire tmp5084;
    wire tmp5085;
    wire tmp5086;
    wire tmp5087;
    wire tmp5088;
    wire tmp5089;
    wire tmp5090;
    wire[254:0] tmp5091;
    wire[255:0] tmp5092;
    wire[256:0] tmp5093;
    wire tmp5094;
    wire tmp5095;
    wire tmp5096;
    wire tmp5097;
    wire tmp5098;
    wire tmp5099;
    wire tmp5100;
    wire tmp5101;
    wire tmp5102;
    wire tmp5103;
    wire[254:0] tmp5104;
    wire[255:0] tmp5105;
    wire[256:0] tmp5106;
    wire tmp5107;
    wire tmp5108;
    wire tmp5109;
    wire tmp5110;
    wire tmp5111;
    wire tmp5112;
    wire tmp5113;
    wire tmp5114;
    wire[254:0] tmp5115;
    wire[255:0] tmp5116;
    wire tmp5117;
    wire[256:0] tmp5118;
    wire tmp5119;
    wire tmp5120;
    wire tmp5121;
    wire tmp5122;
    wire tmp5123;
    wire tmp5124;
    wire tmp5125;
    wire tmp5126;
    wire tmp5127;
    wire tmp5128;
    wire[255:0] tmp5129;
    wire[255:0] tmp5130;
    wire tmp5131;
    wire tmp5132;
    wire tmp5133;
    wire tmp5134;
    wire tmp5135;
    wire tmp5136;
    wire tmp5137;
    wire tmp5138;
    wire tmp5139;
    wire tmp5140;
    wire tmp5141;
    wire tmp5142;
    wire tmp5143;
    wire tmp5144;
    wire tmp5145;
    wire tmp5146;
    wire tmp5147;
    wire tmp5148;
    wire tmp5149;
    wire tmp5150;
    wire tmp5151;
    wire tmp5152;
    wire tmp5153;
    wire[254:0] tmp5154;
    wire[255:0] tmp5155;
    wire tmp5156;
    wire[254:0] tmp5157;
    wire[255:0] tmp5158;
    wire tmp5159;
    wire[256:0] tmp5160;
    wire tmp5161;
    wire tmp5162;
    wire tmp5163;
    wire tmp5164;
    wire tmp5165;
    wire tmp5166;
    wire tmp5167;
    wire tmp5168;
    wire tmp5169;
    wire[254:0] tmp5170;
    wire[255:0] tmp5171;
    wire[256:0] tmp5172;
    wire tmp5173;
    wire tmp5174;
    wire tmp5175;
    wire tmp5176;
    wire tmp5177;
    wire tmp5178;
    wire tmp5179;
    wire tmp5180;
    wire tmp5181;
    wire tmp5182;
    wire[254:0] tmp5183;
    wire[255:0] tmp5184;
    wire[256:0] tmp5185;
    wire tmp5186;
    wire tmp5187;
    wire tmp5188;
    wire tmp5189;
    wire tmp5190;
    wire tmp5191;
    wire tmp5192;
    wire tmp5193;
    wire[254:0] tmp5194;
    wire[255:0] tmp5195;
    wire tmp5196;
    wire[256:0] tmp5197;
    wire tmp5198;
    wire tmp5199;
    wire tmp5200;
    wire tmp5201;
    wire tmp5202;
    wire tmp5203;
    wire tmp5204;
    wire tmp5205;
    wire tmp5206;
    wire tmp5207;
    wire[255:0] tmp5208;
    wire[255:0] tmp5209;
    wire tmp5210;
    wire tmp5211;
    wire[256:0] tmp5212;
    wire tmp5213;
    wire tmp5214;
    wire tmp5215;
    wire tmp5216;
    wire tmp5217;
    wire tmp5218;
    wire tmp5219;
    wire[254:0] tmp5220;
    wire[255:0] tmp5221;
    wire tmp5222;
    wire[254:0] tmp5223;
    wire[255:0] tmp5224;
    wire tmp5225;
    wire[256:0] tmp5226;
    wire tmp5227;
    wire tmp5228;
    wire tmp5229;
    wire tmp5230;
    wire tmp5231;
    wire tmp5232;
    wire tmp5233;
    wire tmp5234;
    wire tmp5235;
    wire[254:0] tmp5236;
    wire[255:0] tmp5237;
    wire[256:0] tmp5238;
    wire tmp5239;
    wire tmp5240;
    wire tmp5241;
    wire tmp5242;
    wire tmp5243;
    wire tmp5244;
    wire tmp5245;
    wire tmp5246;
    wire tmp5247;
    wire tmp5248;
    wire[254:0] tmp5249;
    wire[255:0] tmp5250;
    wire[256:0] tmp5251;
    wire tmp5252;
    wire tmp5253;
    wire tmp5254;
    wire tmp5255;
    wire tmp5256;
    wire tmp5257;
    wire tmp5258;
    wire tmp5259;
    wire[254:0] tmp5260;
    wire[255:0] tmp5261;
    wire tmp5262;
    wire[256:0] tmp5263;
    wire tmp5264;
    wire tmp5265;
    wire tmp5266;
    wire tmp5267;
    wire tmp5268;
    wire tmp5269;
    wire tmp5270;
    wire tmp5271;
    wire tmp5272;
    wire tmp5273;
    wire[255:0] tmp5274;
    wire[255:0] tmp5275;
    wire tmp5276;
    wire tmp5277;
    wire[256:0] tmp5278;
    wire tmp5279;
    wire tmp5280;
    wire tmp5281;
    wire tmp5282;
    wire tmp5283;
    wire tmp5284;
    wire tmp5285;
    wire tmp5286;
    wire[254:0] tmp5287;
    wire[255:0] tmp5288;
    wire tmp5289;
    wire[254:0] tmp5290;
    wire[255:0] tmp5291;
    wire tmp5292;
    wire[256:0] tmp5293;
    wire tmp5294;
    wire tmp5295;
    wire tmp5296;
    wire tmp5297;
    wire tmp5298;
    wire tmp5299;
    wire tmp5300;
    wire tmp5301;
    wire tmp5302;
    wire[254:0] tmp5303;
    wire[255:0] tmp5304;
    wire[256:0] tmp5305;
    wire tmp5306;
    wire tmp5307;
    wire tmp5308;
    wire tmp5309;
    wire tmp5310;
    wire tmp5311;
    wire tmp5312;
    wire tmp5313;
    wire tmp5314;
    wire tmp5315;
    wire[254:0] tmp5316;
    wire[255:0] tmp5317;
    wire[256:0] tmp5318;
    wire tmp5319;
    wire tmp5320;
    wire tmp5321;
    wire tmp5322;
    wire tmp5323;
    wire tmp5324;
    wire tmp5325;
    wire tmp5326;
    wire[254:0] tmp5327;
    wire[255:0] tmp5328;
    wire tmp5329;
    wire[256:0] tmp5330;
    wire tmp5331;
    wire tmp5332;
    wire tmp5333;
    wire tmp5334;
    wire tmp5335;
    wire tmp5336;
    wire tmp5337;
    wire tmp5338;
    wire tmp5339;
    wire tmp5340;
    wire[255:0] tmp5341;
    wire[255:0] tmp5342;
    wire tmp5343;
    wire tmp5344;
    wire[256:0] tmp5345;
    wire tmp5346;
    wire tmp5347;
    wire tmp5348;
    wire tmp5349;
    wire tmp5350;
    wire tmp5351;
    wire tmp5352;
    wire tmp5353;
    wire[254:0] tmp5354;
    wire[255:0] tmp5355;
    wire tmp5356;
    wire[254:0] tmp5357;
    wire[255:0] tmp5358;
    wire tmp5359;
    wire[256:0] tmp5360;
    wire tmp5361;
    wire tmp5362;
    wire tmp5363;
    wire tmp5364;
    wire tmp5365;
    wire tmp5366;
    wire tmp5367;
    wire tmp5368;
    wire tmp5369;
    wire[254:0] tmp5370;
    wire[255:0] tmp5371;
    wire[256:0] tmp5372;
    wire tmp5373;
    wire tmp5374;
    wire tmp5375;
    wire tmp5376;
    wire tmp5377;
    wire tmp5378;
    wire tmp5379;
    wire tmp5380;
    wire tmp5381;
    wire tmp5382;
    wire[254:0] tmp5383;
    wire[255:0] tmp5384;
    wire[256:0] tmp5385;
    wire tmp5386;
    wire tmp5387;
    wire tmp5388;
    wire tmp5389;
    wire tmp5390;
    wire tmp5391;
    wire tmp5392;
    wire tmp5393;
    wire[254:0] tmp5394;
    wire[255:0] tmp5395;
    wire tmp5396;
    wire[256:0] tmp5397;
    wire tmp5398;
    wire tmp5399;
    wire tmp5400;
    wire tmp5401;
    wire tmp5402;
    wire tmp5403;
    wire tmp5404;
    wire tmp5405;
    wire tmp5406;
    wire tmp5407;
    wire[255:0] tmp5408;
    wire[255:0] tmp5409;
    wire tmp5410;
    wire tmp5411;
    wire[256:0] tmp5412;
    wire tmp5413;
    wire tmp5414;
    wire tmp5415;
    wire tmp5416;
    wire tmp5417;
    wire tmp5418;
    wire tmp5419;
    wire tmp5420;
    wire[254:0] tmp5421;
    wire[255:0] tmp5422;
    wire tmp5423;
    wire[254:0] tmp5424;
    wire[255:0] tmp5425;
    wire tmp5426;
    wire[256:0] tmp5427;
    wire tmp5428;
    wire tmp5429;
    wire tmp5430;
    wire tmp5431;
    wire tmp5432;
    wire tmp5433;
    wire tmp5434;
    wire tmp5435;
    wire tmp5436;
    wire[254:0] tmp5437;
    wire[255:0] tmp5438;
    wire[256:0] tmp5439;
    wire tmp5440;
    wire tmp5441;
    wire tmp5442;
    wire tmp5443;
    wire tmp5444;
    wire tmp5445;
    wire tmp5446;
    wire tmp5447;
    wire tmp5448;
    wire tmp5449;
    wire[254:0] tmp5450;
    wire[255:0] tmp5451;
    wire[256:0] tmp5452;
    wire tmp5453;
    wire tmp5454;
    wire tmp5455;
    wire tmp5456;
    wire tmp5457;
    wire tmp5458;
    wire tmp5459;
    wire tmp5460;
    wire[254:0] tmp5461;
    wire[255:0] tmp5462;
    wire tmp5463;
    wire[256:0] tmp5464;
    wire tmp5465;
    wire tmp5466;
    wire tmp5467;
    wire tmp5468;
    wire tmp5469;
    wire tmp5470;
    wire tmp5471;
    wire tmp5472;
    wire tmp5473;
    wire tmp5474;
    wire[255:0] tmp5475;
    wire[255:0] tmp5476;
    wire tmp5477;
    wire tmp5478;
    wire[256:0] tmp5479;
    wire tmp5480;
    wire tmp5481;
    wire tmp5482;
    wire tmp5483;
    wire tmp5484;
    wire tmp5485;
    wire tmp5486;
    wire tmp5487;
    wire[254:0] tmp5488;
    wire[255:0] tmp5489;
    wire tmp5490;
    wire[254:0] tmp5491;
    wire[255:0] tmp5492;
    wire tmp5493;
    wire[256:0] tmp5494;
    wire tmp5495;
    wire tmp5496;
    wire tmp5497;
    wire tmp5498;
    wire tmp5499;
    wire tmp5500;
    wire tmp5501;
    wire tmp5502;
    wire tmp5503;
    wire[254:0] tmp5504;
    wire[255:0] tmp5505;
    wire[256:0] tmp5506;
    wire tmp5507;
    wire tmp5508;
    wire tmp5509;
    wire tmp5510;
    wire tmp5511;
    wire tmp5512;
    wire tmp5513;
    wire tmp5514;
    wire tmp5515;
    wire tmp5516;
    wire[254:0] tmp5517;
    wire[255:0] tmp5518;
    wire[256:0] tmp5519;
    wire tmp5520;
    wire tmp5521;
    wire tmp5522;
    wire tmp5523;
    wire tmp5524;
    wire tmp5525;
    wire tmp5526;
    wire tmp5527;
    wire[254:0] tmp5528;
    wire[255:0] tmp5529;
    wire tmp5530;
    wire[256:0] tmp5531;
    wire tmp5532;
    wire tmp5533;
    wire tmp5534;
    wire tmp5535;
    wire tmp5536;
    wire tmp5537;
    wire tmp5538;
    wire tmp5539;
    wire tmp5540;
    wire tmp5541;
    wire[255:0] tmp5542;
    wire[255:0] tmp5543;
    wire tmp5544;
    wire tmp5545;
    wire[256:0] tmp5546;
    wire tmp5547;
    wire tmp5548;
    wire tmp5549;
    wire tmp5550;
    wire tmp5551;
    wire tmp5552;
    wire tmp5553;
    wire tmp5554;
    wire[254:0] tmp5555;
    wire[255:0] tmp5556;
    wire tmp5557;
    wire[254:0] tmp5558;
    wire[255:0] tmp5559;
    wire tmp5560;
    wire[256:0] tmp5561;
    wire tmp5562;
    wire tmp5563;
    wire tmp5564;
    wire tmp5565;
    wire tmp5566;
    wire tmp5567;
    wire tmp5568;
    wire tmp5569;
    wire tmp5570;
    wire[254:0] tmp5571;
    wire[255:0] tmp5572;
    wire[256:0] tmp5573;
    wire tmp5574;
    wire tmp5575;
    wire tmp5576;
    wire tmp5577;
    wire tmp5578;
    wire tmp5579;
    wire tmp5580;
    wire tmp5581;
    wire tmp5582;
    wire tmp5583;
    wire[254:0] tmp5584;
    wire[255:0] tmp5585;
    wire[256:0] tmp5586;
    wire tmp5587;
    wire tmp5588;
    wire tmp5589;
    wire tmp5590;
    wire tmp5591;
    wire tmp5592;
    wire tmp5593;
    wire tmp5594;
    wire[254:0] tmp5595;
    wire[255:0] tmp5596;
    wire tmp5597;
    wire[256:0] tmp5598;
    wire tmp5599;
    wire tmp5600;
    wire tmp5601;
    wire tmp5602;
    wire tmp5603;
    wire tmp5604;
    wire tmp5605;
    wire tmp5606;
    wire tmp5607;
    wire tmp5608;
    wire[255:0] tmp5609;
    wire[255:0] tmp5610;
    wire tmp5611;
    wire tmp5612;
    wire[256:0] tmp5613;
    wire tmp5614;
    wire tmp5615;
    wire tmp5616;
    wire tmp5617;
    wire tmp5618;
    wire tmp5619;
    wire tmp5620;
    wire tmp5621;
    wire[254:0] tmp5622;
    wire[255:0] tmp5623;
    wire tmp5624;
    wire[254:0] tmp5625;
    wire[255:0] tmp5626;
    wire tmp5627;
    wire[256:0] tmp5628;
    wire tmp5629;
    wire tmp5630;
    wire tmp5631;
    wire tmp5632;
    wire tmp5633;
    wire tmp5634;
    wire tmp5635;
    wire tmp5636;
    wire tmp5637;
    wire[254:0] tmp5638;
    wire[255:0] tmp5639;
    wire[256:0] tmp5640;
    wire tmp5641;
    wire tmp5642;
    wire tmp5643;
    wire tmp5644;
    wire tmp5645;
    wire tmp5646;
    wire tmp5647;
    wire tmp5648;
    wire tmp5649;
    wire tmp5650;
    wire[254:0] tmp5651;
    wire[255:0] tmp5652;
    wire[256:0] tmp5653;
    wire tmp5654;
    wire tmp5655;
    wire tmp5656;
    wire tmp5657;
    wire tmp5658;
    wire tmp5659;
    wire tmp5660;
    wire tmp5661;
    wire[254:0] tmp5662;
    wire[255:0] tmp5663;
    wire tmp5664;
    wire[256:0] tmp5665;
    wire tmp5666;
    wire tmp5667;
    wire tmp5668;
    wire tmp5669;
    wire tmp5670;
    wire tmp5671;
    wire tmp5672;
    wire tmp5673;
    wire tmp5674;
    wire tmp5675;
    wire[255:0] tmp5676;
    wire[255:0] tmp5677;
    wire tmp5678;
    wire tmp5679;
    wire[256:0] tmp5680;
    wire tmp5681;
    wire tmp5682;
    wire tmp5683;
    wire tmp5684;
    wire tmp5685;
    wire tmp5686;
    wire tmp5687;
    wire tmp5688;
    wire tmp5689;
    wire tmp5690;
    wire tmp5691;
    wire tmp5692;
    wire tmp5693;
    wire tmp5694;
    wire tmp5695;
    wire tmp5696;
    wire tmp5697;
    wire tmp5698;
    wire tmp5699;
    wire tmp5700;
    wire tmp5701;
    wire tmp5702;
    wire tmp5703;
    wire tmp5704;
    wire tmp5705;
    wire tmp5706;
    wire tmp5707;
    wire tmp5708;
    wire tmp5709;
    wire tmp5710;
    wire tmp5711;
    wire tmp5712;
    wire tmp5713;
    wire tmp5714;
    wire tmp5715;
    wire tmp5716;
    wire tmp5717;
    wire tmp5718;
    wire tmp5719;
    wire tmp5720;
    wire tmp5721;
    wire tmp5722;
    wire tmp5723;
    wire tmp5724;
    wire tmp5725;
    wire tmp5726;
    wire tmp5727;
    wire tmp5728;
    wire tmp5729;
    wire tmp5730;
    wire tmp5731;
    wire tmp5732;
    wire tmp5733;
    wire tmp5734;
    wire tmp5735;
    wire tmp5736;
    wire tmp5737;
    wire tmp5738;
    wire tmp5739;
    wire tmp5740;
    wire tmp5741;
    wire tmp5742;
    wire tmp5743;
    wire tmp5744;
    wire tmp5745;
    wire tmp5746;
    wire tmp5747;
    wire tmp5748;
    wire tmp5749;
    wire tmp5750;
    wire tmp5751;
    wire tmp5752;
    wire tmp5753;
    wire tmp5754;
    wire tmp5755;
    wire tmp5756;
    wire tmp5757;
    wire tmp5758;
    wire[254:0] tmp5759;
    wire[255:0] tmp5760;
    wire[256:0] tmp5761;
    wire[1:0] tmp5762;
    wire[256:0] tmp5763;
    wire[256:0] tmp5764;
    wire tmp5765;
    wire[1:0] tmp5766;
    wire[257:0] tmp5767;
    wire tmp5768;
    wire tmp5769;
    wire[257:0] tmp5770;
    wire[258:0] tmp5771;
    wire[257:0] tmp5772;
    wire[255:0] tmp5773;
    wire tmp5774;
    wire[254:0] tmp5775;
    wire[255:0] tmp5776;
    wire tmp5777;
    wire[256:0] tmp5778;
    wire tmp5779;
    wire tmp5780;
    wire tmp5781;
    wire tmp5782;
    wire tmp5783;
    wire tmp5784;
    wire tmp5785;
    wire tmp5786;
    wire[255:0] tmp5787;
    wire[256:0] tmp5788;
    wire tmp5789;
    wire[257:0] tmp5790;
    wire tmp5791;
    wire tmp5792;
    wire tmp5793;
    wire tmp5794;
    wire tmp5795;
    wire tmp5796;
    wire tmp5797;
    wire tmp5798;
    wire tmp5799;
    wire tmp5800;
    wire[254:0] tmp5801;
    wire[255:0] tmp5802;
    wire[256:0] tmp5803;
    wire tmp5804;
    wire tmp5805;
    wire tmp5806;
    wire tmp5807;
    wire tmp5808;
    wire tmp5809;
    wire tmp5810;
    wire tmp5811;
    wire tmp5812;
    wire tmp5813;
    wire tmp5814;
    wire tmp5815;
    wire[254:0] tmp5816;
    wire[255:0] tmp5817;
    wire[256:0] tmp5818;
    wire tmp5819;
    wire tmp5820;
    wire tmp5821;
    wire tmp5822;
    wire tmp5823;
    wire tmp5824;
    wire tmp5825;
    wire tmp5826;
    wire tmp5827;
    wire[255:0] tmp5828;
    wire[256:0] tmp5829;
    wire[257:0] tmp5830;
    wire tmp5831;
    wire tmp5832;
    wire tmp5833;
    wire tmp5834;
    wire tmp5835;
    wire tmp5836;
    wire tmp5837;
    wire tmp5838;
    wire tmp5839;
    wire[254:0] tmp5840;
    wire[255:0] tmp5841;
    wire tmp5842;
    wire[256:0] tmp5843;
    wire tmp5844;
    wire tmp5845;
    wire tmp5846;
    wire tmp5847;
    wire tmp5848;
    wire tmp5849;
    wire tmp5850;
    wire tmp5851;
    wire tmp5852;
    wire tmp5853;
    wire[255:0] tmp5854;
    wire[255:0] tmp5855;
    wire tmp5856;
    wire tmp5857;
    wire tmp5858;
    wire tmp5859;
    wire tmp5860;
    wire tmp5861;
    wire tmp5862;
    wire tmp5863;
    wire tmp5864;
    wire tmp5865;
    wire tmp5866;
    wire tmp5867;
    wire tmp5868;
    wire tmp5869;
    wire tmp5870;
    wire tmp5871;
    wire tmp5872;
    wire tmp5873;
    wire tmp5874;
    wire tmp5875;
    wire tmp5876;
    wire tmp5877;
    wire tmp5878;
    wire tmp5879;
    wire tmp5880;
    wire tmp5881;
    wire tmp5882;
    wire tmp5883;
    wire tmp5884;
    wire tmp5885;
    wire tmp5886;
    wire tmp5887;
    wire tmp5888;
    wire tmp5889;
    wire tmp5890;
    wire tmp5891;
    wire tmp5892;
    wire tmp5893;
    wire tmp5894;
    wire tmp5895;
    wire tmp5896;
    wire tmp5897;
    wire tmp5898;
    wire tmp5899;
    wire tmp5900;
    wire tmp5901;
    wire tmp5902;
    wire[254:0] tmp5903;
    wire[255:0] tmp5904;
    wire[256:0] tmp5905;
    wire[1:0] tmp5906;
    wire[256:0] tmp5907;
    wire[256:0] tmp5908;
    wire tmp5909;
    wire[1:0] tmp5910;
    wire[257:0] tmp5911;
    wire tmp5912;
    wire tmp5913;
    wire[257:0] tmp5914;
    wire[258:0] tmp5915;
    wire[257:0] tmp5916;
    wire[255:0] tmp5917;
    wire tmp5918;
    wire[254:0] tmp5919;
    wire[255:0] tmp5920;
    wire tmp5921;
    wire[256:0] tmp5922;
    wire tmp5923;
    wire tmp5924;
    wire tmp5925;
    wire tmp5926;
    wire tmp5927;
    wire tmp5928;
    wire tmp5929;
    wire tmp5930;
    wire[255:0] tmp5931;
    wire[256:0] tmp5932;
    wire tmp5933;
    wire[257:0] tmp5934;
    wire tmp5935;
    wire tmp5936;
    wire tmp5937;
    wire tmp5938;
    wire tmp5939;
    wire tmp5940;
    wire tmp5941;
    wire tmp5942;
    wire tmp5943;
    wire tmp5944;
    wire[254:0] tmp5945;
    wire[255:0] tmp5946;
    wire[256:0] tmp5947;
    wire tmp5948;
    wire tmp5949;
    wire tmp5950;
    wire tmp5951;
    wire tmp5952;
    wire tmp5953;
    wire tmp5954;
    wire tmp5955;
    wire tmp5956;
    wire tmp5957;
    wire tmp5958;
    wire tmp5959;
    wire[254:0] tmp5960;
    wire[255:0] tmp5961;
    wire[256:0] tmp5962;
    wire tmp5963;
    wire tmp5964;
    wire tmp5965;
    wire tmp5966;
    wire tmp5967;
    wire tmp5968;
    wire tmp5969;
    wire tmp5970;
    wire tmp5971;
    wire[255:0] tmp5972;
    wire[256:0] tmp5973;
    wire[257:0] tmp5974;
    wire tmp5975;
    wire tmp5976;
    wire tmp5977;
    wire tmp5978;
    wire tmp5979;
    wire tmp5980;
    wire tmp5981;
    wire tmp5982;
    wire tmp5983;
    wire[254:0] tmp5984;
    wire[255:0] tmp5985;
    wire tmp5986;
    wire[256:0] tmp5987;
    wire tmp5988;
    wire tmp5989;
    wire tmp5990;
    wire tmp5991;
    wire tmp5992;
    wire tmp5993;
    wire tmp5994;
    wire tmp5995;
    wire tmp5996;
    wire tmp5997;
    wire[255:0] tmp5998;
    wire[255:0] tmp5999;
    wire tmp6000;
    wire tmp6001;
    wire tmp6002;
    wire tmp6003;
    wire tmp6004;
    wire tmp6005;
    wire tmp6006;
    wire tmp6007;
    wire tmp6008;
    wire tmp6009;
    wire tmp6010;
    wire tmp6011;
    wire tmp6012;
    wire tmp6013;
    wire tmp6014;
    wire tmp6015;
    wire tmp6016;
    wire tmp6017;
    wire tmp6018;
    wire tmp6019;
    wire tmp6020;
    wire tmp6021;
    wire tmp6022;
    wire tmp6023;
    wire tmp6024;
    wire tmp6025;
    wire tmp6026;
    wire tmp6027;
    wire tmp6028;
    wire tmp6029;
    wire tmp6030;
    wire tmp6031;
    wire tmp6032;
    wire tmp6033;
    wire tmp6034;
    wire tmp6035;
    wire tmp6036;
    wire tmp6037;
    wire tmp6038;
    wire tmp6039;
    wire tmp6040;
    wire tmp6041;
    wire tmp6042;
    wire tmp6043;
    wire tmp6044;
    wire tmp6045;
    wire tmp6046;
    wire[254:0] tmp6047;
    wire[255:0] tmp6048;
    wire[256:0] tmp6049;
    wire[1:0] tmp6050;
    wire[256:0] tmp6051;
    wire[256:0] tmp6052;
    wire tmp6053;
    wire[1:0] tmp6054;
    wire[257:0] tmp6055;
    wire tmp6056;
    wire tmp6057;
    wire[257:0] tmp6058;
    wire[258:0] tmp6059;
    wire[257:0] tmp6060;
    wire[255:0] tmp6061;
    wire tmp6062;
    wire[254:0] tmp6063;
    wire[255:0] tmp6064;
    wire tmp6065;
    wire[256:0] tmp6066;
    wire tmp6067;
    wire tmp6068;
    wire tmp6069;
    wire tmp6070;
    wire tmp6071;
    wire tmp6072;
    wire tmp6073;
    wire tmp6074;
    wire[255:0] tmp6075;
    wire[256:0] tmp6076;
    wire tmp6077;
    wire[257:0] tmp6078;
    wire tmp6079;
    wire tmp6080;
    wire tmp6081;
    wire tmp6082;
    wire tmp6083;
    wire tmp6084;
    wire tmp6085;
    wire tmp6086;
    wire tmp6087;
    wire tmp6088;
    wire[254:0] tmp6089;
    wire[255:0] tmp6090;
    wire[256:0] tmp6091;
    wire tmp6092;
    wire tmp6093;
    wire tmp6094;
    wire tmp6095;
    wire tmp6096;
    wire tmp6097;
    wire tmp6098;
    wire tmp6099;
    wire tmp6100;
    wire tmp6101;
    wire tmp6102;
    wire tmp6103;
    wire[254:0] tmp6104;
    wire[255:0] tmp6105;
    wire[256:0] tmp6106;
    wire tmp6107;
    wire tmp6108;
    wire tmp6109;
    wire tmp6110;
    wire tmp6111;
    wire tmp6112;
    wire tmp6113;
    wire tmp6114;
    wire tmp6115;
    wire[255:0] tmp6116;
    wire[256:0] tmp6117;
    wire[257:0] tmp6118;
    wire tmp6119;
    wire tmp6120;
    wire tmp6121;
    wire tmp6122;
    wire tmp6123;
    wire tmp6124;
    wire tmp6125;
    wire tmp6126;
    wire tmp6127;
    wire[254:0] tmp6128;
    wire[255:0] tmp6129;
    wire tmp6130;
    wire[256:0] tmp6131;
    wire tmp6132;
    wire tmp6133;
    wire tmp6134;
    wire tmp6135;
    wire tmp6136;
    wire tmp6137;
    wire tmp6138;
    wire tmp6139;
    wire tmp6140;
    wire tmp6141;
    wire[255:0] tmp6142;
    wire[255:0] tmp6143;
    wire tmp6144;
    wire tmp6145;
    wire tmp6146;
    wire tmp6147;
    wire tmp6148;
    wire tmp6149;
    wire tmp6150;
    wire tmp6151;
    wire tmp6152;
    wire tmp6153;
    wire tmp6154;
    wire tmp6155;
    wire tmp6156;
    wire tmp6157;
    wire tmp6158;
    wire tmp6159;
    wire tmp6160;
    wire tmp6161;
    wire tmp6162;
    wire tmp6163;
    wire tmp6164;
    wire tmp6165;
    wire tmp6166;
    wire tmp6167;
    wire tmp6168;
    wire tmp6169;
    wire tmp6170;
    wire tmp6171;
    wire tmp6172;
    wire tmp6173;
    wire tmp6174;
    wire tmp6175;
    wire tmp6176;
    wire tmp6177;
    wire tmp6178;
    wire tmp6179;
    wire tmp6180;
    wire tmp6181;
    wire tmp6182;
    wire tmp6183;
    wire tmp6184;
    wire tmp6185;
    wire tmp6186;
    wire tmp6187;
    wire tmp6188;
    wire tmp6189;
    wire tmp6190;
    wire[254:0] tmp6191;
    wire[255:0] tmp6192;
    wire[256:0] tmp6193;
    wire[1:0] tmp6194;
    wire[256:0] tmp6195;
    wire[256:0] tmp6196;
    wire tmp6197;
    wire[1:0] tmp6198;
    wire[257:0] tmp6199;
    wire tmp6200;
    wire tmp6201;
    wire[257:0] tmp6202;
    wire[258:0] tmp6203;
    wire[257:0] tmp6204;
    wire[255:0] tmp6205;
    wire tmp6206;
    wire[254:0] tmp6207;
    wire[255:0] tmp6208;
    wire tmp6209;
    wire[256:0] tmp6210;
    wire tmp6211;
    wire tmp6212;
    wire tmp6213;
    wire tmp6214;
    wire tmp6215;
    wire tmp6216;
    wire tmp6217;
    wire tmp6218;
    wire[255:0] tmp6219;
    wire[256:0] tmp6220;
    wire tmp6221;
    wire[257:0] tmp6222;
    wire tmp6223;
    wire tmp6224;
    wire tmp6225;
    wire tmp6226;
    wire tmp6227;
    wire tmp6228;
    wire tmp6229;
    wire tmp6230;
    wire tmp6231;
    wire tmp6232;
    wire[254:0] tmp6233;
    wire[255:0] tmp6234;
    wire[256:0] tmp6235;
    wire tmp6236;
    wire tmp6237;
    wire tmp6238;
    wire tmp6239;
    wire tmp6240;
    wire tmp6241;
    wire tmp6242;
    wire tmp6243;
    wire tmp6244;
    wire tmp6245;
    wire tmp6246;
    wire tmp6247;
    wire[254:0] tmp6248;
    wire[255:0] tmp6249;
    wire[256:0] tmp6250;
    wire tmp6251;
    wire tmp6252;
    wire tmp6253;
    wire tmp6254;
    wire tmp6255;
    wire tmp6256;
    wire tmp6257;
    wire tmp6258;
    wire tmp6259;
    wire[255:0] tmp6260;
    wire[256:0] tmp6261;
    wire[257:0] tmp6262;
    wire tmp6263;
    wire tmp6264;
    wire tmp6265;
    wire tmp6266;
    wire tmp6267;
    wire tmp6268;
    wire tmp6269;
    wire tmp6270;
    wire tmp6271;
    wire[254:0] tmp6272;
    wire[255:0] tmp6273;
    wire tmp6274;
    wire[256:0] tmp6275;
    wire tmp6276;
    wire tmp6277;
    wire tmp6278;
    wire tmp6279;
    wire tmp6280;
    wire tmp6281;
    wire tmp6282;
    wire tmp6283;
    wire tmp6284;
    wire tmp6285;
    wire[255:0] tmp6286;
    wire[255:0] tmp6287;
    wire tmp6288;
    wire tmp6289;
    wire tmp6290;
    wire tmp6291;
    wire tmp6292;
    wire tmp6293;
    wire tmp6294;
    wire tmp6295;
    wire tmp6296;
    wire tmp6297;
    wire tmp6298;
    wire tmp6299;
    wire tmp6300;
    wire tmp6301;
    wire tmp6302;
    wire tmp6303;
    wire tmp6304;
    wire tmp6305;
    wire tmp6306;
    wire tmp6307;
    wire tmp6308;
    wire tmp6309;
    wire tmp6310;
    wire tmp6311;
    wire tmp6312;
    wire tmp6313;
    wire tmp6314;
    wire tmp6315;
    wire tmp6316;
    wire tmp6317;
    wire tmp6318;
    wire tmp6319;
    wire tmp6320;
    wire tmp6321;
    wire tmp6322;
    wire tmp6323;
    wire tmp6324;
    wire tmp6325;
    wire tmp6326;
    wire tmp6327;
    wire tmp6328;
    wire tmp6329;
    wire tmp6330;
    wire tmp6331;
    wire tmp6332;
    wire tmp6333;
    wire tmp6334;
    wire tmp6335;
    wire tmp6336;
    wire tmp6337;
    wire tmp6338;
    wire tmp6339;
    wire tmp6340;
    wire tmp6341;
    wire tmp6342;
    wire tmp6343;
    wire tmp6344;
    wire tmp6345;
    wire tmp6346;
    wire tmp6347;
    wire tmp6348;
    wire tmp6349;
    wire tmp6350;
    wire tmp6351;
    wire tmp6352;
    wire tmp6353;
    wire tmp6354;
    wire tmp6355;
    wire tmp6356;
    wire tmp6357;
    wire tmp6358;
    wire tmp6359;
    wire tmp6360;
    wire tmp6361;
    wire tmp6362;
    wire tmp6363;
    wire tmp6364;
    wire tmp6365;
    wire tmp6366;
    wire tmp6367;
    wire tmp6368;
    wire tmp6369;
    wire tmp6370;
    wire tmp6371;
    wire tmp6372;
    wire tmp6373;
    wire tmp6374;
    wire tmp6375;
    wire tmp6376;
    wire tmp6377;
    wire tmp6378;
    wire tmp6379;
    wire tmp6380;
    wire tmp6381;
    wire tmp6382;
    wire tmp6383;
    wire tmp6384;
    wire tmp6385;
    wire tmp6386;
    wire tmp6387;
    wire tmp6388;
    wire tmp6389;
    wire tmp6390;
    wire tmp6391;
    wire tmp6392;
    wire tmp6393;
    wire tmp6394;
    wire tmp6395;
    wire tmp6396;
    wire tmp6397;
    wire tmp6398;
    wire tmp6399;
    wire tmp6400;
    wire tmp6401;
    wire tmp6402;
    wire[254:0] tmp6403;
    wire[255:0] tmp6404;
    wire[256:0] tmp6405;
    wire tmp6406;
    wire tmp6407;
    wire tmp6408;
    wire tmp6409;
    wire tmp6410;
    wire tmp6411;
    wire tmp6412;
    wire tmp6413;
    wire[254:0] tmp6414;
    wire[255:0] tmp6415;
    wire[256:0] tmp6416;
    wire[1:0] tmp6417;
    wire[256:0] tmp6418;
    wire[256:0] tmp6419;
    wire tmp6420;
    wire[256:0] tmp6421;
    wire[256:0] tmp6422;
    wire tmp6423;
    wire tmp6424;
    wire[254:0] tmp6425;
    wire[255:0] tmp6426;
    wire[256:0] tmp6427;
    wire tmp6428;
    wire tmp6429;
    wire tmp6430;
    wire tmp6431;
    wire tmp6432;
    wire tmp6433;
    wire tmp6434;
    wire tmp6435;
    wire[254:0] tmp6436;
    wire[255:0] tmp6437;
    wire[256:0] tmp6438;
    wire[1:0] tmp6439;
    wire[256:0] tmp6440;
    wire[256:0] tmp6441;
    wire tmp6442;
    wire[256:0] tmp6443;
    wire[256:0] tmp6444;
    wire tmp6445;
    wire tmp6446;
    wire[257:0] tmp6447;
    wire tmp6448;
    wire tmp6449;
    wire tmp6450;
    wire tmp6451;
    wire tmp6452;
    wire tmp6453;
    wire tmp6454;
    wire tmp6455;
    wire tmp6456;
    wire[254:0] tmp6457;
    wire[255:0] tmp6458;
    wire[256:0] tmp6459;
    wire tmp6460;
    wire tmp6461;
    wire tmp6462;
    wire tmp6463;
    wire tmp6464;
    wire tmp6465;
    wire tmp6466;
    wire tmp6467;
    wire[254:0] tmp6468;
    wire[255:0] tmp6469;
    wire[256:0] tmp6470;
    wire[1:0] tmp6471;
    wire[256:0] tmp6472;
    wire[256:0] tmp6473;
    wire tmp6474;
    wire[256:0] tmp6475;
    wire[256:0] tmp6476;
    wire tmp6477;
    wire tmp6478;
    wire[254:0] tmp6479;
    wire[255:0] tmp6480;
    wire[256:0] tmp6481;
    wire tmp6482;
    wire tmp6483;
    wire tmp6484;
    wire tmp6485;
    wire tmp6486;
    wire tmp6487;
    wire tmp6488;
    wire tmp6489;
    wire[254:0] tmp6490;
    wire[255:0] tmp6491;
    wire[256:0] tmp6492;
    wire[1:0] tmp6493;
    wire[256:0] tmp6494;
    wire[256:0] tmp6495;
    wire tmp6496;
    wire[256:0] tmp6497;
    wire[256:0] tmp6498;
    wire tmp6499;
    wire tmp6500;
    wire[257:0] tmp6501;
    wire tmp6502;
    wire tmp6503;
    wire tmp6504;
    wire tmp6505;
    wire tmp6506;
    wire tmp6507;
    wire tmp6508;
    wire tmp6509;
    wire tmp6510;
    wire tmp6511;
    wire[254:0] tmp6512;
    wire[255:0] tmp6513;
    wire[256:0] tmp6514;
    wire tmp6515;
    wire tmp6516;
    wire tmp6517;
    wire tmp6518;
    wire tmp6519;
    wire tmp6520;
    wire tmp6521;
    wire tmp6522;
    wire[254:0] tmp6523;
    wire[255:0] tmp6524;
    wire[256:0] tmp6525;
    wire[1:0] tmp6526;
    wire[256:0] tmp6527;
    wire[256:0] tmp6528;
    wire tmp6529;
    wire[256:0] tmp6530;
    wire[256:0] tmp6531;
    wire tmp6532;
    wire tmp6533;
    wire[254:0] tmp6534;
    wire[255:0] tmp6535;
    wire[256:0] tmp6536;
    wire tmp6537;
    wire tmp6538;
    wire tmp6539;
    wire tmp6540;
    wire tmp6541;
    wire tmp6542;
    wire tmp6543;
    wire tmp6544;
    wire[254:0] tmp6545;
    wire[255:0] tmp6546;
    wire[256:0] tmp6547;
    wire[1:0] tmp6548;
    wire[256:0] tmp6549;
    wire[256:0] tmp6550;
    wire tmp6551;
    wire[256:0] tmp6552;
    wire[256:0] tmp6553;
    wire tmp6554;
    wire tmp6555;
    wire[257:0] tmp6556;
    wire tmp6557;
    wire tmp6558;
    wire tmp6559;
    wire tmp6560;
    wire tmp6561;
    wire tmp6562;
    wire tmp6563;
    wire tmp6564;
    wire tmp6565;
    wire tmp6566;
    wire[254:0] tmp6567;
    wire[255:0] tmp6568;
    wire[256:0] tmp6569;
    wire tmp6570;
    wire tmp6571;
    wire tmp6572;
    wire tmp6573;
    wire tmp6574;
    wire tmp6575;
    wire tmp6576;
    wire tmp6577;
    wire[254:0] tmp6578;
    wire[255:0] tmp6579;
    wire[256:0] tmp6580;
    wire[1:0] tmp6581;
    wire[256:0] tmp6582;
    wire[256:0] tmp6583;
    wire tmp6584;
    wire[256:0] tmp6585;
    wire[256:0] tmp6586;
    wire tmp6587;
    wire tmp6588;
    wire[254:0] tmp6589;
    wire[255:0] tmp6590;
    wire[256:0] tmp6591;
    wire tmp6592;
    wire tmp6593;
    wire tmp6594;
    wire tmp6595;
    wire tmp6596;
    wire tmp6597;
    wire tmp6598;
    wire tmp6599;
    wire[254:0] tmp6600;
    wire[255:0] tmp6601;
    wire[256:0] tmp6602;
    wire[1:0] tmp6603;
    wire[256:0] tmp6604;
    wire[256:0] tmp6605;
    wire tmp6606;
    wire[256:0] tmp6607;
    wire[256:0] tmp6608;
    wire tmp6609;
    wire tmp6610;
    wire[257:0] tmp6611;
    wire tmp6612;
    wire tmp6613;
    wire tmp6614;
    wire tmp6615;
    wire tmp6616;
    wire tmp6617;
    wire tmp6618;
    wire tmp6619;
    wire tmp6620;
    wire tmp6621;
    wire tmp6622;
    wire tmp6623;
    wire tmp6624;
    wire tmp6625;
    wire tmp6626;
    wire tmp6627;
    wire tmp6628;
    wire tmp6629;
    wire tmp6630;
    wire tmp6631;
    wire tmp6632;
    wire tmp6633;
    wire tmp6634;
    wire tmp6635;
    wire tmp6636;
    wire tmp6637;
    wire tmp6638;
    wire tmp6639;
    wire tmp6640;
    wire tmp6641;
    wire tmp6642;
    wire tmp6643;
    wire tmp6644;
    wire tmp6645;
    wire tmp6646;
    wire tmp6647;
    wire tmp6648;
    wire tmp6649;
    wire tmp6650;
    wire tmp6651;
    wire tmp6652;
    wire tmp6653;
    wire tmp6654;
    wire tmp6655;
    wire tmp6656;
    wire tmp6657;
    wire tmp6658;
    wire tmp6659;
    wire tmp6660;
    wire tmp6661;
    wire tmp6662;
    wire tmp6663;
    wire tmp6664;
    wire tmp6665;
    wire tmp6666;
    wire tmp6667;
    wire tmp6668;
    wire tmp6669;
    wire tmp6670;
    wire tmp6671;
    wire tmp6672;
    wire tmp6673;
    wire tmp6674;
    wire tmp6675;
    wire tmp6676;
    wire tmp6677;
    wire tmp6678;
    wire tmp6679;
    wire tmp6680;
    wire tmp6681;
    wire tmp6682;
    wire tmp6683;
    wire tmp6684;
    wire tmp6685;
    wire tmp6686;
    wire tmp6687;
    wire tmp6688;
    wire tmp6689;
    wire tmp6690;
    wire tmp6691;
    wire tmp6692;
    wire tmp6693;
    wire tmp6694;
    wire tmp6695;
    wire tmp6696;
    wire tmp6697;
    wire tmp6698;
    wire tmp6699;
    wire tmp6700;
    wire tmp6701;
    wire tmp6702;
    wire tmp6703;
    wire tmp6704;
    wire tmp6705;
    wire tmp6706;
    wire tmp6707;
    wire tmp6708;
    wire tmp6709;
    wire tmp6710;
    wire tmp6711;
    wire tmp6712;
    wire tmp6713;
    wire tmp6714;
    wire tmp6715;
    wire tmp6716;
    wire tmp6717;
    wire tmp6718;
    wire tmp6719;
    wire tmp6720;
    wire tmp6721;
    wire tmp6722;
    wire tmp6723;
    wire tmp6724;
    wire tmp6725;
    wire tmp6726;
    wire tmp6727;
    wire tmp6728;
    wire tmp6729;
    wire tmp6730;
    wire tmp6731;
    wire tmp6732;
    wire tmp6733;
    wire tmp6734;
    wire tmp6735;
    wire tmp6736;
    wire tmp6737;
    wire tmp6738;
    wire tmp6739;
    wire tmp6740;
    wire tmp6741;
    wire tmp6742;
    wire tmp6743;
    wire tmp6744;
    wire tmp6745;
    wire tmp6746;
    wire tmp6747;
    wire tmp6748;
    wire tmp6749;
    wire tmp6750;
    wire tmp6751;
    wire tmp6752;
    wire tmp6753;
    wire tmp6754;
    wire tmp6755;
    wire tmp6756;
    wire tmp6757;
    wire tmp6758;
    wire tmp6759;
    wire tmp6760;
    wire tmp6761;
    wire[254:0] tmp6762;
    wire[255:0] tmp6763;
    wire[256:0] tmp6764;
    wire tmp6765;
    wire tmp6766;
    wire tmp6767;
    wire tmp6768;
    wire tmp6769;
    wire tmp6770;
    wire tmp6771;
    wire tmp6772;
    wire[254:0] tmp6773;
    wire[255:0] tmp6774;
    wire[256:0] tmp6775;
    wire[1:0] tmp6776;
    wire[256:0] tmp6777;
    wire[256:0] tmp6778;
    wire tmp6779;
    wire[256:0] tmp6780;
    wire[256:0] tmp6781;
    wire[255:0] tmp6782;
    wire tmp6783;
    wire tmp6784;
    wire[256:0] tmp6785;
    wire tmp6786;
    wire tmp6787;
    wire[254:0] tmp6788;
    wire[255:0] tmp6789;
    wire[256:0] tmp6790;
    wire tmp6791;
    wire tmp6792;
    wire tmp6793;
    wire tmp6794;
    wire tmp6795;
    wire tmp6796;
    wire tmp6797;
    wire tmp6798;
    wire[254:0] tmp6799;
    wire[255:0] tmp6800;
    wire[256:0] tmp6801;
    wire[1:0] tmp6802;
    wire[256:0] tmp6803;
    wire[256:0] tmp6804;
    wire tmp6805;
    wire[256:0] tmp6806;
    wire[256:0] tmp6807;
    wire tmp6808;
    wire tmp6809;
    wire[257:0] tmp6810;
    wire tmp6811;
    wire tmp6812;
    wire tmp6813;
    wire tmp6814;
    wire tmp6815;
    wire tmp6816;
    wire tmp6817;
    wire tmp6818;
    wire tmp6819;
    wire tmp6820;
    wire tmp6821;
    wire tmp6822;
    wire[254:0] tmp6823;
    wire[255:0] tmp6824;
    wire[256:0] tmp6825;
    wire tmp6826;
    wire tmp6827;
    wire tmp6828;
    wire tmp6829;
    wire tmp6830;
    wire tmp6831;
    wire tmp6832;
    wire tmp6833;
    wire[254:0] tmp6834;
    wire[255:0] tmp6835;
    wire[256:0] tmp6836;
    wire[1:0] tmp6837;
    wire[256:0] tmp6838;
    wire[256:0] tmp6839;
    wire tmp6840;
    wire[256:0] tmp6841;
    wire[256:0] tmp6842;
    wire[255:0] tmp6843;
    wire tmp6844;
    wire tmp6845;
    wire[256:0] tmp6846;
    wire tmp6847;
    wire tmp6848;
    wire[254:0] tmp6849;
    wire[255:0] tmp6850;
    wire[256:0] tmp6851;
    wire tmp6852;
    wire tmp6853;
    wire tmp6854;
    wire tmp6855;
    wire tmp6856;
    wire tmp6857;
    wire tmp6858;
    wire tmp6859;
    wire[254:0] tmp6860;
    wire[255:0] tmp6861;
    wire[256:0] tmp6862;
    wire[1:0] tmp6863;
    wire[256:0] tmp6864;
    wire[256:0] tmp6865;
    wire tmp6866;
    wire[256:0] tmp6867;
    wire[256:0] tmp6868;
    wire tmp6869;
    wire tmp6870;
    wire[257:0] tmp6871;
    wire tmp6872;
    wire tmp6873;
    wire tmp6874;
    wire tmp6875;
    wire tmp6876;
    wire tmp6877;
    wire tmp6878;
    wire tmp6879;
    wire tmp6880;
    wire tmp6881;
    wire tmp6882;
    wire tmp6883;
    wire[254:0] tmp6884;
    wire[255:0] tmp6885;
    wire[256:0] tmp6886;
    wire tmp6887;
    wire tmp6888;
    wire tmp6889;
    wire tmp6890;
    wire tmp6891;
    wire tmp6892;
    wire tmp6893;
    wire tmp6894;
    wire[254:0] tmp6895;
    wire[255:0] tmp6896;
    wire[256:0] tmp6897;
    wire[1:0] tmp6898;
    wire[256:0] tmp6899;
    wire[256:0] tmp6900;
    wire tmp6901;
    wire[256:0] tmp6902;
    wire[256:0] tmp6903;
    wire[255:0] tmp6904;
    wire tmp6905;
    wire tmp6906;
    wire[256:0] tmp6907;
    wire tmp6908;
    wire tmp6909;
    wire[254:0] tmp6910;
    wire[255:0] tmp6911;
    wire[256:0] tmp6912;
    wire tmp6913;
    wire tmp6914;
    wire tmp6915;
    wire tmp6916;
    wire tmp6917;
    wire tmp6918;
    wire tmp6919;
    wire tmp6920;
    wire[254:0] tmp6921;
    wire[255:0] tmp6922;
    wire[256:0] tmp6923;
    wire[1:0] tmp6924;
    wire[256:0] tmp6925;
    wire[256:0] tmp6926;
    wire tmp6927;
    wire[256:0] tmp6928;
    wire[256:0] tmp6929;
    wire tmp6930;
    wire tmp6931;
    wire[257:0] tmp6932;
    wire tmp6933;
    wire tmp6934;
    wire tmp6935;
    wire tmp6936;
    wire tmp6937;
    wire tmp6938;
    wire tmp6939;
    wire tmp6940;
    wire tmp6941;
    wire tmp6942;
    wire tmp6943;
    wire tmp6944;
    wire[254:0] tmp6945;
    wire[255:0] tmp6946;
    wire[256:0] tmp6947;
    wire tmp6948;
    wire tmp6949;
    wire tmp6950;
    wire tmp6951;
    wire tmp6952;
    wire tmp6953;
    wire tmp6954;
    wire tmp6955;
    wire[254:0] tmp6956;
    wire[255:0] tmp6957;
    wire[256:0] tmp6958;
    wire[1:0] tmp6959;
    wire[256:0] tmp6960;
    wire[256:0] tmp6961;
    wire tmp6962;
    wire[256:0] tmp6963;
    wire[256:0] tmp6964;
    wire[255:0] tmp6965;
    wire tmp6966;
    wire tmp6967;
    wire[256:0] tmp6968;
    wire tmp6969;
    wire tmp6970;
    wire[254:0] tmp6971;
    wire[255:0] tmp6972;
    wire[256:0] tmp6973;
    wire tmp6974;
    wire tmp6975;
    wire tmp6976;
    wire tmp6977;
    wire tmp6978;
    wire tmp6979;
    wire tmp6980;
    wire tmp6981;
    wire[254:0] tmp6982;
    wire[255:0] tmp6983;
    wire[256:0] tmp6984;
    wire[1:0] tmp6985;
    wire[256:0] tmp6986;
    wire[256:0] tmp6987;
    wire tmp6988;
    wire[256:0] tmp6989;
    wire[256:0] tmp6990;
    wire tmp6991;
    wire tmp6992;
    wire[257:0] tmp6993;
    wire tmp6994;
    wire tmp6995;
    wire tmp6996;
    wire tmp6997;
    wire tmp6998;
    wire tmp6999;
    wire tmp7000;
    wire tmp7001;
    wire tmp7002;
    wire tmp7003;
    wire tmp7004;
    wire tmp7005;
    wire tmp7006;
    wire tmp7007;
    wire tmp7008;
    wire tmp7009;
    wire tmp7010;
    wire tmp7011;
    wire tmp7012;
    wire tmp7013;
    wire tmp7014;
    wire tmp7015;
    wire tmp7016;
    wire tmp7017;
    wire tmp7018;
    wire tmp7019;
    wire tmp7020;
    wire tmp7021;
    wire tmp7022;
    wire tmp7023;
    wire tmp7024;
    wire tmp7025;
    wire tmp7026;
    wire tmp7027;
    wire tmp7028;
    wire tmp7029;
    wire tmp7030;
    wire tmp7031;
    wire tmp7032;
    wire tmp7033;
    wire tmp7034;
    wire tmp7035;
    wire[254:0] tmp7036;
    wire tmp7037;
    wire tmp7038;
    wire[255:0] tmp7039;
    wire tmp7040;
    wire tmp7041;
    wire tmp7042;
    wire tmp7043;
    wire tmp7044;
    wire tmp7045;
    wire tmp7046;
    wire tmp7047;
    wire tmp7048;
    wire tmp7049;
    wire tmp7050;
    wire tmp7051;
    wire tmp7052;
    wire tmp7053;
    wire tmp7054;
    wire tmp7055;
    wire tmp7056;
    wire[254:0] tmp7057;
    wire tmp7058;
    wire tmp7059;
    wire[255:0] tmp7060;
    wire tmp7061;
    wire tmp7062;
    wire tmp7063;
    wire tmp7064;
    wire tmp7065;
    wire tmp7066;
    wire tmp7067;
    wire tmp7068;
    wire tmp7069;
    wire tmp7070;
    wire tmp7071;
    wire tmp7072;
    wire tmp7073;
    wire tmp7074;
    wire tmp7075;
    wire tmp7076;
    wire tmp7077;
    wire[254:0] tmp7078;
    wire tmp7079;
    wire tmp7080;
    wire[255:0] tmp7081;
    wire tmp7082;
    wire tmp7083;
    wire tmp7084;
    wire tmp7085;
    wire tmp7086;
    wire tmp7087;
    wire tmp7088;
    wire tmp7089;
    wire tmp7090;
    wire tmp7091;
    wire tmp7092;
    wire tmp7093;
    wire tmp7094;
    wire tmp7095;
    wire tmp7096;
    wire tmp7097;
    wire tmp7098;
    wire[254:0] tmp7099;
    wire tmp7100;
    wire tmp7101;
    wire[255:0] tmp7102;
    wire tmp7103;
    wire tmp7104;
    wire tmp7105;
    wire tmp7106;
    wire tmp7107;
    wire tmp7108;
    wire tmp7109;
    wire tmp7110;
    wire tmp7111;
    wire tmp7112;
    wire tmp7113;
    wire tmp7114;
    wire tmp7115;
    wire tmp7116;
    wire tmp7117;
    wire tmp7118;
    wire tmp7119;
    wire[254:0] tmp7120;
    wire[255:0] tmp7121;
    wire tmp7122;
    wire[254:0] tmp7123;
    wire[255:0] tmp7124;
    wire tmp7125;
    wire[256:0] tmp7126;
    wire tmp7127;
    wire tmp7128;
    wire tmp7129;
    wire tmp7130;
    wire tmp7131;
    wire tmp7132;
    wire tmp7133;
    wire tmp7134;
    wire tmp7135;
    wire[254:0] tmp7136;
    wire[255:0] tmp7137;
    wire[256:0] tmp7138;
    wire tmp7139;
    wire tmp7140;
    wire tmp7141;
    wire tmp7142;
    wire tmp7143;
    wire tmp7144;
    wire tmp7145;
    wire tmp7146;
    wire tmp7147;
    wire tmp7148;
    wire[254:0] tmp7149;
    wire[255:0] tmp7150;
    wire[256:0] tmp7151;
    wire tmp7152;
    wire tmp7153;
    wire tmp7154;
    wire tmp7155;
    wire tmp7156;
    wire tmp7157;
    wire tmp7158;
    wire tmp7159;
    wire[254:0] tmp7160;
    wire[255:0] tmp7161;
    wire tmp7162;
    wire[256:0] tmp7163;
    wire tmp7164;
    wire tmp7165;
    wire tmp7166;
    wire tmp7167;
    wire tmp7168;
    wire tmp7169;
    wire tmp7170;
    wire tmp7171;
    wire tmp7172;
    wire tmp7173;
    wire[255:0] tmp7174;
    wire[255:0] tmp7175;
    wire tmp7176;
    wire tmp7177;
    wire tmp7178;
    wire tmp7179;
    wire tmp7180;
    wire tmp7181;
    wire tmp7182;
    wire tmp7183;
    wire tmp7184;
    wire tmp7185;
    wire tmp7186;
    wire tmp7187;
    wire tmp7188;
    wire tmp7189;
    wire tmp7190;
    wire tmp7191;
    wire tmp7192;
    wire tmp7193;
    wire[254:0] tmp7194;
    wire[255:0] tmp7195;
    wire tmp7196;
    wire[254:0] tmp7197;
    wire[255:0] tmp7198;
    wire tmp7199;
    wire[256:0] tmp7200;
    wire tmp7201;
    wire tmp7202;
    wire tmp7203;
    wire tmp7204;
    wire tmp7205;
    wire tmp7206;
    wire tmp7207;
    wire tmp7208;
    wire tmp7209;
    wire[254:0] tmp7210;
    wire[255:0] tmp7211;
    wire[256:0] tmp7212;
    wire tmp7213;
    wire tmp7214;
    wire tmp7215;
    wire tmp7216;
    wire tmp7217;
    wire tmp7218;
    wire tmp7219;
    wire tmp7220;
    wire tmp7221;
    wire tmp7222;
    wire[254:0] tmp7223;
    wire[255:0] tmp7224;
    wire[256:0] tmp7225;
    wire tmp7226;
    wire tmp7227;
    wire tmp7228;
    wire tmp7229;
    wire tmp7230;
    wire tmp7231;
    wire tmp7232;
    wire tmp7233;
    wire[254:0] tmp7234;
    wire[255:0] tmp7235;
    wire tmp7236;
    wire[256:0] tmp7237;
    wire tmp7238;
    wire tmp7239;
    wire tmp7240;
    wire tmp7241;
    wire tmp7242;
    wire tmp7243;
    wire tmp7244;
    wire tmp7245;
    wire tmp7246;
    wire tmp7247;
    wire[255:0] tmp7248;
    wire[255:0] tmp7249;
    wire tmp7250;
    wire tmp7251;
    wire tmp7252;
    wire tmp7253;
    wire tmp7254;
    wire tmp7255;
    wire tmp7256;
    wire tmp7257;
    wire tmp7258;
    wire tmp7259;
    wire tmp7260;
    wire tmp7261;
    wire tmp7262;
    wire tmp7263;
    wire tmp7264;
    wire tmp7265;
    wire tmp7266;
    wire tmp7267;
    wire[254:0] tmp7268;
    wire[255:0] tmp7269;
    wire tmp7270;
    wire[254:0] tmp7271;
    wire[255:0] tmp7272;
    wire tmp7273;
    wire[256:0] tmp7274;
    wire tmp7275;
    wire tmp7276;
    wire tmp7277;
    wire tmp7278;
    wire tmp7279;
    wire tmp7280;
    wire tmp7281;
    wire tmp7282;
    wire tmp7283;
    wire[254:0] tmp7284;
    wire[255:0] tmp7285;
    wire[256:0] tmp7286;
    wire tmp7287;
    wire tmp7288;
    wire tmp7289;
    wire tmp7290;
    wire tmp7291;
    wire tmp7292;
    wire tmp7293;
    wire tmp7294;
    wire tmp7295;
    wire tmp7296;
    wire[254:0] tmp7297;
    wire[255:0] tmp7298;
    wire[256:0] tmp7299;
    wire tmp7300;
    wire tmp7301;
    wire tmp7302;
    wire tmp7303;
    wire tmp7304;
    wire tmp7305;
    wire tmp7306;
    wire tmp7307;
    wire[254:0] tmp7308;
    wire[255:0] tmp7309;
    wire tmp7310;
    wire[256:0] tmp7311;
    wire tmp7312;
    wire tmp7313;
    wire tmp7314;
    wire tmp7315;
    wire tmp7316;
    wire tmp7317;
    wire tmp7318;
    wire tmp7319;
    wire tmp7320;
    wire tmp7321;
    wire[255:0] tmp7322;
    wire[255:0] tmp7323;
    wire tmp7324;
    wire tmp7325;
    wire tmp7326;
    wire tmp7327;
    wire tmp7328;
    wire tmp7329;
    wire tmp7330;
    wire tmp7331;
    wire tmp7332;
    wire tmp7333;
    wire tmp7334;
    wire tmp7335;
    wire tmp7336;
    wire tmp7337;
    wire tmp7338;
    wire tmp7339;
    wire tmp7340;
    wire tmp7341;
    wire[254:0] tmp7342;
    wire[255:0] tmp7343;
    wire tmp7344;
    wire[254:0] tmp7345;
    wire[255:0] tmp7346;
    wire tmp7347;
    wire[256:0] tmp7348;
    wire tmp7349;
    wire tmp7350;
    wire tmp7351;
    wire tmp7352;
    wire tmp7353;
    wire tmp7354;
    wire tmp7355;
    wire tmp7356;
    wire tmp7357;
    wire[254:0] tmp7358;
    wire[255:0] tmp7359;
    wire[256:0] tmp7360;
    wire tmp7361;
    wire tmp7362;
    wire tmp7363;
    wire tmp7364;
    wire tmp7365;
    wire tmp7366;
    wire tmp7367;
    wire tmp7368;
    wire tmp7369;
    wire tmp7370;
    wire[254:0] tmp7371;
    wire[255:0] tmp7372;
    wire[256:0] tmp7373;
    wire tmp7374;
    wire tmp7375;
    wire tmp7376;
    wire tmp7377;
    wire tmp7378;
    wire tmp7379;
    wire tmp7380;
    wire tmp7381;
    wire[254:0] tmp7382;
    wire[255:0] tmp7383;
    wire tmp7384;
    wire[256:0] tmp7385;
    wire tmp7386;
    wire tmp7387;
    wire tmp7388;
    wire tmp7389;
    wire tmp7390;
    wire tmp7391;
    wire tmp7392;
    wire tmp7393;
    wire tmp7394;
    wire tmp7395;
    wire[255:0] tmp7396;
    wire[255:0] tmp7397;
    wire tmp7398;
    wire tmp7399;
    wire tmp7400;
    wire tmp7401;
    wire tmp7402;
    wire tmp7403;
    wire tmp7404;
    wire tmp7405;
    wire tmp7406;
    wire tmp7407;
    wire tmp7408;
    wire tmp7409;
    wire tmp7410;
    wire tmp7411;
    wire tmp7412;
    wire tmp7413;
    wire tmp7414;
    wire tmp7415;
    wire tmp7416;
    wire tmp7417;
    wire tmp7418;
    wire tmp7419;
    wire tmp7420;
    wire tmp7421;
    wire tmp7422;
    wire tmp7423;
    wire tmp7424;
    wire tmp7425;
    wire tmp7426;
    wire tmp7427;
    wire tmp7428;
    wire tmp7429;
    wire tmp7430;
    wire tmp7431;
    wire tmp7432;
    wire tmp7433;
    wire tmp7434;
    wire tmp7435;
    wire tmp7436;
    wire tmp7437;
    wire tmp7438;
    wire tmp7439;
    wire tmp7440;
    wire tmp7441;
    wire tmp7442;
    wire tmp7443;
    wire tmp7444;
    wire tmp7445;
    wire tmp7446;
    wire tmp7447;
    wire tmp7448;
    wire tmp7449;
    wire tmp7450;
    wire tmp7451;
    wire tmp7452;
    wire tmp7453;
    wire tmp7454;
    wire tmp7455;
    wire tmp7456;
    wire tmp7457;
    wire tmp7458;
    wire tmp7459;
    wire tmp7460;
    wire tmp7461;
    wire tmp7462;
    wire tmp7463;
    wire tmp7464;
    wire tmp7465;
    wire tmp7466;
    wire tmp7467;
    wire tmp7468;
    wire tmp7469;
    wire tmp7470;
    wire tmp7471;
    wire tmp7472;
    wire tmp7473;
    wire tmp7474;
    wire tmp7475;
    wire tmp7476;
    wire tmp7477;
    wire[255:0] tmp7478;
    wire[255:0] tmp7479;
    wire[255:0] tmp7480;
    wire[255:0] tmp7481;
    wire[255:0] tmp7482;
    wire[255:0] tmp7483;
    wire[255:0] tmp7484;
    wire[255:0] tmp7485;
    wire[255:0] tmp7486;
    wire[255:0] tmp7487;
    wire[255:0] tmp7488;
    wire[255:0] tmp7489;
    wire[255:0] tmp7490;
    wire[255:0] tmp7491;
    wire[255:0] tmp7492;
    wire[255:0] tmp7493;
    wire[255:0] tmp7494;
    wire[255:0] tmp7495;
    wire[255:0] tmp7496;
    wire[255:0] tmp7497;
    wire[255:0] tmp7498;
    wire[255:0] tmp7499;
    wire[255:0] tmp7500;
    wire[255:0] tmp7501;
    wire[255:0] tmp7502;
    wire[255:0] tmp7503;
    wire[255:0] tmp7504;
    wire[255:0] tmp7505;
    wire[255:0] tmp7506;
    wire[255:0] tmp7507;
    wire[255:0] tmp7508;
    wire[255:0] tmp7509;
    wire[255:0] tmp7510;
    wire[255:0] tmp7511;
    wire[255:0] tmp7512;
    wire[255:0] tmp7513;
    wire[255:0] tmp7514;
    wire[255:0] tmp7515;
    wire[255:0] tmp7516;
    wire[255:0] tmp7517;
    wire[255:0] tmp7518;
    wire[255:0] tmp7519;
    wire[255:0] tmp7520;
    wire[255:0] tmp7521;
    wire[255:0] tmp7522;
    wire[255:0] tmp7523;
    wire[255:0] tmp7524;
    wire[255:0] tmp7525;
    wire[255:0] tmp7526;
    wire[255:0] tmp7527;
    wire[255:0] tmp7528;
    wire[255:0] tmp7529;
    wire[255:0] tmp7530;
    wire[255:0] tmp7531;
    wire[255:0] tmp7532;
    wire[255:0] tmp7533;
    wire[255:0] tmp7534;
    wire[255:0] tmp7535;
    wire[255:0] tmp7536;
    wire[255:0] tmp7537;
    wire[255:0] tmp7538;
    wire[255:0] tmp7539;
    wire[255:0] tmp7540;
    wire[255:0] tmp7541;
    wire[255:0] tmp7542;
    wire[255:0] tmp7543;
    wire[255:0] tmp7544;
    wire[255:0] tmp7545;
    wire[255:0] tmp7546;
    wire[255:0] tmp7547;
    wire[255:0] tmp7548;
    wire[255:0] tmp7549;
    wire[255:0] tmp7550;
    wire[255:0] tmp7551;
    wire[255:0] tmp7552;
    wire[255:0] tmp7553;
    wire[255:0] tmp7554;
    wire[255:0] tmp7555;
    wire[255:0] tmp7556;
    wire[255:0] tmp7557;
    wire[255:0] tmp7558;
    wire[255:0] tmp7559;
    wire[255:0] tmp7560;
    wire[255:0] tmp7561;
    wire[255:0] tmp7562;
    wire[255:0] tmp7563;
    wire[255:0] tmp7564;
    wire[255:0] tmp7565;
    wire[255:0] tmp7566;
    wire[255:0] tmp7567;
    wire[255:0] tmp7568;
    wire[255:0] tmp7569;
    wire[255:0] tmp7570;
    wire[255:0] tmp7571;
    wire[255:0] tmp7572;
    wire[255:0] tmp7573;
    wire[255:0] tmp7574;
    wire[255:0] tmp7575;
    wire[255:0] tmp7576;
    wire[255:0] tmp7577;
    wire[255:0] tmp7578;
    wire[255:0] tmp7579;
    wire[255:0] tmp7580;
    wire[255:0] tmp7581;
    wire[255:0] tmp7582;
    wire[255:0] tmp7583;
    wire[255:0] tmp7584;
    wire[255:0] tmp7585;
    wire[255:0] tmp7586;
    wire[255:0] tmp7587;
    wire[255:0] tmp7588;
    wire[255:0] tmp7589;
    wire[255:0] tmp7590;
    wire[255:0] tmp7591;
    wire[255:0] tmp7592;
    wire[255:0] tmp7593;
    wire[255:0] tmp7594;
    wire[255:0] tmp7595;
    wire[255:0] tmp7596;
    wire[255:0] tmp7597;
    wire[255:0] tmp7598;
    wire[255:0] tmp7599;
    wire[255:0] tmp7600;
    wire[255:0] tmp7601;
    wire[255:0] tmp7602;
    wire[255:0] tmp7603;
    wire[255:0] tmp7604;
    wire[255:0] tmp7605;
    wire[255:0] tmp7606;
    wire[255:0] tmp7607;
    wire[255:0] tmp7608;
    wire[255:0] tmp7609;
    wire[255:0] tmp7610;
    wire[255:0] tmp7611;
    wire[255:0] tmp7612;
    wire[255:0] tmp7613;
    wire[255:0] tmp7614;
    wire[255:0] tmp7615;
    wire[255:0] tmp7616;
    wire[255:0] tmp7617;
    wire tmp7618;
    wire tmp7619;
    wire tmp7620;
    wire tmp7621;
    wire tmp7622;
    wire tmp7623;
    wire tmp7624;
    wire tmp7625;
    wire tmp7626;
    wire tmp7627;
    wire tmp7628;
    wire tmp7629;
    wire tmp7630;
    wire tmp7631;
    wire tmp7632;
    wire tmp7633;
    wire[2:0] tmp7634;
    wire[3:0] tmp7635;
    wire[3:0] tmp7636;
    wire[3:0] tmp7637;
    wire[3:0] tmp7638;
    wire[3:0] tmp7639;
    wire[3:0] tmp7640;
    wire[3:0] tmp7641;
    wire[3:0] tmp7642;
    wire[3:0] tmp7643;
    wire[3:0] tmp7644;
    wire[3:0] tmp7645;
    wire[3:0] tmp7646;
    wire[3:0] tmp7647;
    wire[3:0] tmp7648;
    wire[3:0] tmp7649;
    wire[3:0] tmp7650;
    wire tmp7651;
    wire tmp7652;
    wire tmp7653;
    wire tmp7654;
    wire tmp7655;
    wire[254:0] tmp7656;
    wire[255:0] tmp7657;
    wire[255:0] tmp7658;
    wire[255:0] tmp7659;
    wire[254:0] tmp7660;
    wire[255:0] tmp7661;
    wire[255:0] tmp7662;
    wire[255:0] tmp7663;
    wire[254:0] tmp7664;
    wire[255:0] tmp7665;
    wire[255:0] tmp7666;
    wire[255:0] tmp7667;
    wire[254:0] tmp7668;
    wire[255:0] tmp7669;
    wire[255:0] tmp7670;
    wire[255:0] tmp7671;
    wire[254:0] tmp7672;
    wire[255:0] tmp7673;
    wire[255:0] tmp7674;
    wire[255:0] tmp7675;
    wire[254:0] tmp7676;
    wire[255:0] tmp7677;
    wire[255:0] tmp7678;
    wire[255:0] tmp7679;
    wire[254:0] tmp7680;
    wire[255:0] tmp7681;
    wire[255:0] tmp7682;
    wire[255:0] tmp7683;
    wire[254:0] tmp7684;
    wire[255:0] tmp7685;
    wire[255:0] tmp7686;
    wire[255:0] tmp7687;
    wire[1:0] tmp7689;
    wire[2:0] tmp7690;
    wire tmp7691;
    wire tmp7692;
    wire[2:0] tmp7693;
    wire tmp7694;
    wire tmp7695;
    wire tmp7696;
    wire[2:0] tmp7697;
    wire tmp7698;
    wire tmp7699;
    wire tmp7700;
    wire[3:0] tmp7701;
    wire tmp7702;
    wire tmp7703;
    wire tmp7704;
    wire tmp7705;
    wire tmp7706;
    wire tmp7707;
    wire tmp7708;
    wire tmp7709;
    wire tmp7710;
    wire tmp7711;
    wire[3:0] tmp7712;
    wire tmp7713;
    wire tmp7714;
    wire tmp7715;
    wire[3:0] tmp7716;
    wire tmp7717;
    wire tmp7718;
    wire tmp7719;
    wire tmp7720;
    wire tmp7721;
    wire tmp7722;
    wire[3:0] tmp7723;
    wire tmp7724;
    wire tmp7725;
    wire[1:0] tmp7726;
    wire[2:0] tmp7727;
    wire tmp7728;
    wire tmp7729;
    wire[1:0] tmp7730;
    wire[2:0] tmp7731;
    wire tmp7732;
    wire tmp7733;
    wire tmp7734;
    wire tmp7735;
    wire tmp7736;
    wire tmp7737;
    wire tmp7738;
    wire tmp7739;
    wire[2:0] tmp7740;
    wire tmp7741;
    wire tmp7742;
    wire tmp7743;
    wire tmp7744;
    wire tmp7745;
    wire tmp7746;
    wire tmp7747;
    wire tmp7748;
    wire tmp7749;
    wire tmp7750;
    wire tmp7751;
    wire[2:0] tmp7752;
    wire tmp7753;
    wire tmp7754;
    wire tmp7755;
    wire tmp7756;
    wire tmp7757;
    wire tmp7758;
    wire[2:0] tmp7759;
    wire tmp7760;
    wire tmp7761;
    wire tmp7762;
    wire tmp7763;
    wire tmp7764;
    wire tmp7765;
    wire tmp7766;
    wire tmp7767;
    wire[1:0] tmp7768;
    wire[2:0] tmp7769;
    wire[2:0] tmp7770;
    wire[2:0] tmp7771;
    wire[2:0] tmp7772;
    wire[2:0] tmp7773;
    wire[2:0] tmp7774;
    wire[3:0] tmp7775;
    wire[3:0] tmp7776;
    wire[2:0] tmp7777;
    wire[3:0] tmp7778;
    wire[3:0] tmp7779;
    wire[2:0] tmp7780;

    // Combinational
    assign _ver_out_tmp_0 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_1 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_2 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_3 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_4 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_5 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_6 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_7 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_8 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_9 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_10 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_11 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_12 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_13 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_14 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_15 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_16 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_17 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_18 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_19 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_20 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_21 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_22 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_23 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_24 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_25 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_26 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_27 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_28 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_29 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_30 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_31 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_32 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_33 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_34 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_35 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_36 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_37 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_38 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_39 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_40 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_41 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_42 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_43 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_44 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_45 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_46 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_47 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_48 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_49 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_50 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_51 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_52 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_53 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_54 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_55 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_56 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_57 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_58 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_59 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_60 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_61 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_62 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_63 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_64 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_65 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_66 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_67 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_68 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_69 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_70 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_71 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_72 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_73 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_74 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_75 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_76 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_77 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_78 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_79 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_80 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_81 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_82 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_83 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_84 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_85 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_86 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_87 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_88 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_89 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_90 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign _ver_out_tmp_91 = 57896044618658097711785492504343953926634992332820282019728792003956564819968;
    assign const_0_1 = 1;
    assign const_1_1 = 1;
    assign const_2_0 = 0;
    assign const_3_0 = 0;
    assign const_4_0 = 0;
    assign const_5_4 = 4;
    assign const_6_0 = 0;
    assign const_7_2 = 2;
    assign const_8_1 = 1;
    assign const_9_0 = 0;
    assign const_10_0 = 0;
    assign const_11_0 = 0;
    assign const_12_0 = 0;
    assign const_13_1 = 1;
    assign const_14_0 = 0;
    assign const_15_1 = 1;
    assign const_16_0 = 0;
    assign const_17_0 = 0;
    assign const_18_0 = 0;
    assign const_19_0 = 0;
    assign const_20_15 = 15;
    assign const_21_1 = 1;
    assign const_22_0 = 0;
    assign const_23_2 = 2;
    assign const_24_0 = 0;
    assign const_25_3 = 3;
    assign const_26_0 = 0;
    assign const_27_0 = 0;
    assign const_28_0 = 0;
    assign const_29_0 = 0;
    assign const_30_0 = 0;
    assign const_31_0 = 0;
    assign const_32_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_34_0 = 0;
    assign const_35_0 = 0;
    assign const_36_0 = 0;
    assign const_37_0 = 0;
    assign const_38_0 = 0;
    assign const_39_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_41_0 = 0;
    assign const_42_0 = 0;
    assign const_43_0 = 0;
    assign const_44_0 = 0;
    assign const_45_0 = 0;
    assign const_46_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_48_0 = 0;
    assign const_49_0 = 0;
    assign const_50_0 = 0;
    assign const_51_0 = 0;
    assign const_52_0 = 0;
    assign const_53_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_55_6 = 6;
    assign const_56_0 = 0;
    assign const_57_7 = 7;
    assign const_58_0 = 0;
    assign const_59_4 = 4;
    assign const_60_0 = 0;
    assign const_61_5 = 5;
    assign const_62_0 = 0;
    assign const_63_0 = 0;
    assign const_64_0 = 0;
    assign const_65_0 = 0;
    assign const_66_0 = 0;
    assign const_67_0 = 0;
    assign const_68_0 = 0;
    assign const_69_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_71_0 = 0;
    assign const_72_0 = 0;
    assign const_73_0 = 0;
    assign const_74_0 = 0;
    assign const_75_0 = 0;
    assign const_76_0 = 0;
    assign const_77_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_79_0 = 0;
    assign const_80_0 = 0;
    assign const_81_0 = 0;
    assign const_82_0 = 0;
    assign const_83_0 = 0;
    assign const_84_0 = 0;
    assign const_85_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_87_0 = 0;
    assign const_88_0 = 0;
    assign const_89_0 = 0;
    assign const_90_0 = 0;
    assign const_91_0 = 0;
    assign const_92_0 = 0;
    assign const_93_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_95_8 = 8;
    assign const_97_0 = 0;
    assign const_98_0 = 0;
    assign const_99_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_100_0 = 0;
    assign const_102_0 = 0;
    assign const_103_0 = 0;
    assign const_104_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_105_0 = 0;
    assign const_107_0 = 0;
    assign const_108_0 = 0;
    assign const_109_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_110_0 = 0;
    assign const_112_0 = 0;
    assign const_113_0 = 0;
    assign const_114_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_115_0 = 0;
    assign const_116_2 = 2;
    assign const_117_0 = 0;
    assign const_118_0 = 0;
    assign const_119_0 = 0;
    assign const_120_0 = 0;
    assign const_121_15 = 15;
    assign const_122_1 = 1;
    assign const_123_0 = 0;
    assign const_124_2 = 2;
    assign const_125_0 = 0;
    assign const_126_3 = 3;
    assign const_127_0 = 0;
    assign const_128_0 = 0;
    assign const_129_0 = 0;
    assign const_130_0 = 0;
    assign const_131_0 = 0;
    assign const_132_0 = 0;
    assign const_133_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_135_0 = 0;
    assign const_136_0 = 0;
    assign const_137_0 = 0;
    assign const_138_0 = 0;
    assign const_139_0 = 0;
    assign const_140_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_142_0 = 0;
    assign const_143_0 = 0;
    assign const_144_0 = 0;
    assign const_145_0 = 0;
    assign const_146_0 = 0;
    assign const_147_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_149_0 = 0;
    assign const_150_0 = 0;
    assign const_151_0 = 0;
    assign const_152_0 = 0;
    assign const_153_0 = 0;
    assign const_154_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_156_6 = 6;
    assign const_157_0 = 0;
    assign const_158_7 = 7;
    assign const_159_0 = 0;
    assign const_160_4 = 4;
    assign const_161_0 = 0;
    assign const_162_5 = 5;
    assign const_163_0 = 0;
    assign const_164_0 = 0;
    assign const_165_0 = 0;
    assign const_166_0 = 0;
    assign const_167_0 = 0;
    assign const_168_0 = 0;
    assign const_169_0 = 0;
    assign const_170_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_172_0 = 0;
    assign const_173_0 = 0;
    assign const_174_0 = 0;
    assign const_175_0 = 0;
    assign const_176_0 = 0;
    assign const_177_0 = 0;
    assign const_178_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_180_0 = 0;
    assign const_181_0 = 0;
    assign const_182_0 = 0;
    assign const_183_0 = 0;
    assign const_184_0 = 0;
    assign const_185_0 = 0;
    assign const_186_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_188_0 = 0;
    assign const_189_0 = 0;
    assign const_190_0 = 0;
    assign const_191_0 = 0;
    assign const_192_0 = 0;
    assign const_193_0 = 0;
    assign const_194_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_196_8 = 8;
    assign const_198_0 = 0;
    assign const_199_0 = 0;
    assign const_200_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_201_0 = 0;
    assign const_203_0 = 0;
    assign const_204_0 = 0;
    assign const_205_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_206_0 = 0;
    assign const_208_0 = 0;
    assign const_209_0 = 0;
    assign const_210_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_211_0 = 0;
    assign const_213_0 = 0;
    assign const_214_0 = 0;
    assign const_215_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_216_0 = 0;
    assign const_217_3 = 3;
    assign const_218_0 = 0;
    assign const_219_0 = 0;
    assign const_220_0 = 0;
    assign const_221_0 = 0;
    assign const_222_0 = 0;
    assign const_223_0 = 0;
    assign const_224_0 = 0;
    assign const_225_0 = 0;
    assign const_226_0 = 0;
    assign const_227_0 = 0;
    assign const_228_0 = 0;
    assign const_229_0 = 0;
    assign const_230_0 = 0;
    assign const_231_0 = 0;
    assign const_232_0 = 0;
    assign const_233_0 = 0;
    assign const_234_0 = 0;
    assign const_235_0 = 0;
    assign const_236_0 = 0;
    assign const_237_0 = 0;
    assign const_238_0 = 0;
    assign const_239_0 = 0;
    assign const_240_0 = 0;
    assign const_242_0 = 0;
    assign const_243_0 = 0;
    assign const_244_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_245_0 = 0;
    assign const_247_0 = 0;
    assign const_248_0 = 0;
    assign const_249_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_250_0 = 0;
    assign const_252_0 = 0;
    assign const_253_0 = 0;
    assign const_254_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_255_0 = 0;
    assign const_257_0 = 0;
    assign const_258_0 = 0;
    assign const_259_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_260_0 = 0;
    assign const_262_0 = 0;
    assign const_263_0 = 0;
    assign const_264_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_265_0 = 0;
    assign const_267_0 = 0;
    assign const_268_0 = 0;
    assign const_269_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_270_0 = 0;
    assign const_272_0 = 0;
    assign const_273_0 = 0;
    assign const_274_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_275_0 = 0;
    assign const_277_0 = 0;
    assign const_278_0 = 0;
    assign const_279_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_280_0 = 0;
    assign const_281_0 = 0;
    assign const_282_0 = 0;
    assign const_283_0 = 0;
    assign const_284_0 = 0;
    assign const_285_0 = 0;
    assign const_286_0 = 0;
    assign const_287_0 = 0;
    assign const_288_0 = 0;
    assign const_289_0 = 0;
    assign const_290_0 = 0;
    assign const_291_15 = 15;
    assign const_292_0 = 0;
    assign const_293_0 = 0;
    assign const_294_0 = 0;
    assign const_295_8 = 8;
    assign const_296_0 = 0;
    assign const_298_0 = 0;
    assign const_299_0 = 0;
    assign const_300_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_301_0 = 0;
    assign const_303_0 = 0;
    assign const_304_0 = 0;
    assign const_305_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_306_0 = 0;
    assign const_308_0 = 0;
    assign const_309_0 = 0;
    assign const_310_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_311_0 = 0;
    assign const_313_0 = 0;
    assign const_314_0 = 0;
    assign const_315_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_316_0 = 0;
    assign const_317_1 = 1;
    assign const_318_0 = 0;
    assign const_319_0 = 0;
    assign const_320_0 = 0;
    assign const_321_0 = 0;
    assign const_322_0 = 0;
    assign const_323_0 = 0;
    assign const_324_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_326_0 = 0;
    assign const_327_0 = 0;
    assign const_328_0 = 0;
    assign const_329_0 = 0;
    assign const_330_0 = 0;
    assign const_331_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_333_0 = 0;
    assign const_334_0 = 0;
    assign const_335_0 = 0;
    assign const_336_0 = 0;
    assign const_337_0 = 0;
    assign const_338_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_340_0 = 0;
    assign const_341_0 = 0;
    assign const_342_0 = 0;
    assign const_343_0 = 0;
    assign const_344_0 = 0;
    assign const_345_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_347_4 = 4;
    assign const_348_0 = 0;
    assign const_350_0 = 0;
    assign const_351_0 = 0;
    assign const_352_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_353_0 = 0;
    assign const_354_0 = 0;
    assign const_355_0 = 0;
    assign const_356_0 = 0;
    assign const_357_0 = 0;
    assign const_358_0 = 0;
    assign const_359_0 = 0;
    assign const_360_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_363_0 = 0;
    assign const_364_0 = 0;
    assign const_365_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_366_0 = 0;
    assign const_367_0 = 0;
    assign const_368_0 = 0;
    assign const_369_0 = 0;
    assign const_370_0 = 0;
    assign const_371_0 = 0;
    assign const_372_0 = 0;
    assign const_373_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_376_0 = 0;
    assign const_377_0 = 0;
    assign const_378_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_379_0 = 0;
    assign const_380_0 = 0;
    assign const_381_0 = 0;
    assign const_382_0 = 0;
    assign const_383_0 = 0;
    assign const_384_0 = 0;
    assign const_385_0 = 0;
    assign const_386_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_389_0 = 0;
    assign const_390_0 = 0;
    assign const_391_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_392_0 = 0;
    assign const_393_0 = 0;
    assign const_394_0 = 0;
    assign const_395_0 = 0;
    assign const_396_0 = 0;
    assign const_397_0 = 0;
    assign const_398_0 = 0;
    assign const_399_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_401_6 = 6;
    assign const_402_0 = 0;
    assign const_403_0 = 0;
    assign const_404_0 = 0;
    assign const_405_0 = 0;
    assign const_406_0 = 0;
    assign const_407_0 = 0;
    assign const_408_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_410_0 = 0;
    assign const_411_0 = 0;
    assign const_412_0 = 0;
    assign const_413_0 = 0;
    assign const_414_0 = 0;
    assign const_415_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_417_0 = 0;
    assign const_418_0 = 0;
    assign const_419_0 = 0;
    assign const_420_0 = 0;
    assign const_421_0 = 0;
    assign const_422_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_424_0 = 0;
    assign const_425_0 = 0;
    assign const_426_0 = 0;
    assign const_427_0 = 0;
    assign const_428_0 = 0;
    assign const_429_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_431_2 = 2;
    assign const_432_0 = 0;
    assign const_433_0 = 0;
    assign const_434_0 = 0;
    assign const_435_0 = 0;
    assign const_436_0 = 0;
    assign const_437_0 = 0;
    assign const_438_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_440_0 = 0;
    assign const_441_0 = 0;
    assign const_442_0 = 0;
    assign const_443_0 = 0;
    assign const_444_0 = 0;
    assign const_445_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_447_0 = 0;
    assign const_448_0 = 0;
    assign const_449_0 = 0;
    assign const_450_0 = 0;
    assign const_451_0 = 0;
    assign const_452_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_454_0 = 0;
    assign const_455_0 = 0;
    assign const_456_0 = 0;
    assign const_457_0 = 0;
    assign const_458_0 = 0;
    assign const_459_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_461_0 = 0;
    assign const_462_0 = 0;
    assign const_463_0 = 0;
    assign const_464_0 = 0;
    assign const_465_0 = 0;
    assign const_466_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_468_0 = 0;
    assign const_469_0 = 0;
    assign const_470_0 = 0;
    assign const_471_0 = 0;
    assign const_472_0 = 0;
    assign const_473_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_475_0 = 0;
    assign const_476_0 = 0;
    assign const_477_0 = 0;
    assign const_478_0 = 0;
    assign const_479_0 = 0;
    assign const_480_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_482_0 = 0;
    assign const_483_0 = 0;
    assign const_484_0 = 0;
    assign const_485_0 = 0;
    assign const_486_0 = 0;
    assign const_487_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_489_0 = 0;
    assign const_490_0 = 0;
    assign const_491_0 = 0;
    assign const_492_0 = 0;
    assign const_493_0 = 0;
    assign const_494_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_496_0 = 0;
    assign const_497_0 = 0;
    assign const_498_0 = 0;
    assign const_499_0 = 0;
    assign const_500_0 = 0;
    assign const_501_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_503_0 = 0;
    assign const_504_0 = 0;
    assign const_505_0 = 0;
    assign const_506_0 = 0;
    assign const_507_0 = 0;
    assign const_508_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_510_0 = 0;
    assign const_511_0 = 0;
    assign const_512_0 = 0;
    assign const_513_0 = 0;
    assign const_514_0 = 0;
    assign const_515_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_517_5 = 5;
    assign const_518_1 = 1;
    assign const_520_0 = 0;
    assign const_521_0 = 0;
    assign const_522_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_523_0 = 0;
    assign const_524_0 = 0;
    assign const_525_0 = 0;
    assign const_526_0 = 0;
    assign const_527_0 = 0;
    assign const_528_0 = 0;
    assign const_529_0 = 0;
    assign const_530_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_533_0 = 0;
    assign const_534_0 = 0;
    assign const_535_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_536_0 = 0;
    assign const_537_0 = 0;
    assign const_538_0 = 0;
    assign const_539_0 = 0;
    assign const_540_0 = 0;
    assign const_541_0 = 0;
    assign const_542_0 = 0;
    assign const_543_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_546_0 = 0;
    assign const_547_0 = 0;
    assign const_548_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_549_0 = 0;
    assign const_550_0 = 0;
    assign const_551_0 = 0;
    assign const_552_0 = 0;
    assign const_553_0 = 0;
    assign const_554_0 = 0;
    assign const_555_0 = 0;
    assign const_556_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_559_0 = 0;
    assign const_560_0 = 0;
    assign const_561_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_562_0 = 0;
    assign const_563_0 = 0;
    assign const_564_0 = 0;
    assign const_565_0 = 0;
    assign const_566_0 = 0;
    assign const_567_0 = 0;
    assign const_568_0 = 0;
    assign const_569_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_571_0 = 0;
    assign const_572_0 = 0;
    assign const_573_0 = 0;
    assign const_574_0 = 0;
    assign const_575_0 = 0;
    assign const_577_0 = 0;
    assign const_578_0 = 0;
    assign const_579_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_580_0 = 0;
    assign const_581_0 = 0;
    assign const_582_0 = 0;
    assign const_584_0 = 0;
    assign const_585_0 = 0;
    assign const_586_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_587_0 = 0;
    assign const_588_0 = 0;
    assign const_589_0 = 0;
    assign const_591_0 = 0;
    assign const_592_0 = 0;
    assign const_593_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_594_0 = 0;
    assign const_595_0 = 0;
    assign const_596_0 = 0;
    assign const_598_0 = 0;
    assign const_599_0 = 0;
    assign const_600_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_601_0 = 0;
    assign const_602_0 = 0;
    assign const_603_0 = 0;
    assign const_605_0 = 0;
    assign const_606_0 = 0;
    assign const_607_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_608_0 = 0;
    assign const_609_0 = 0;
    assign const_610_0 = 0;
    assign const_612_0 = 0;
    assign const_613_0 = 0;
    assign const_614_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_615_0 = 0;
    assign const_616_0 = 0;
    assign const_617_0 = 0;
    assign const_619_0 = 0;
    assign const_620_0 = 0;
    assign const_621_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_622_0 = 0;
    assign const_623_0 = 0;
    assign const_624_0 = 0;
    assign const_626_0 = 0;
    assign const_627_0 = 0;
    assign const_628_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_629_0 = 0;
    assign const_630_0 = 0;
    assign const_631_6 = 6;
    assign const_632_1 = 1;
    assign const_633_0 = 0;
    assign const_635_0 = 0;
    assign const_636_0 = 0;
    assign const_637_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_638_0 = 0;
    assign const_639_0 = 0;
    assign const_640_0 = 0;
    assign const_642_0 = 0;
    assign const_643_0 = 0;
    assign const_644_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_645_0 = 0;
    assign const_646_0 = 0;
    assign const_647_0 = 0;
    assign const_649_0 = 0;
    assign const_650_0 = 0;
    assign const_651_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_652_0 = 0;
    assign const_653_0 = 0;
    assign const_654_0 = 0;
    assign const_656_0 = 0;
    assign const_657_0 = 0;
    assign const_658_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_659_0 = 0;
    assign const_660_0 = 0;
    assign const_661_0 = 0;
    assign const_663_0 = 0;
    assign const_664_0 = 0;
    assign const_665_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_666_0 = 0;
    assign const_667_0 = 0;
    assign const_668_0 = 0;
    assign const_670_0 = 0;
    assign const_671_0 = 0;
    assign const_672_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_673_0 = 0;
    assign const_674_0 = 0;
    assign const_675_0 = 0;
    assign const_677_0 = 0;
    assign const_678_0 = 0;
    assign const_679_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_680_0 = 0;
    assign const_681_0 = 0;
    assign const_682_0 = 0;
    assign const_684_0 = 0;
    assign const_685_0 = 0;
    assign const_686_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_687_0 = 0;
    assign const_688_0 = 0;
    assign const_689_3 = 3;
    assign const_690_1 = 1;
    assign const_691_0 = 0;
    assign const_692_0 = 0;
    assign const_693_0 = 0;
    assign const_694_0 = 0;
    assign const_695_0 = 0;
    assign const_696_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_698_0 = 0;
    assign const_699_0 = 0;
    assign const_700_0 = 0;
    assign const_701_0 = 0;
    assign const_702_0 = 0;
    assign const_703_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_705_0 = 0;
    assign const_706_0 = 0;
    assign const_707_0 = 0;
    assign const_708_0 = 0;
    assign const_709_0 = 0;
    assign const_710_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_712_0 = 0;
    assign const_713_0 = 0;
    assign const_714_0 = 0;
    assign const_715_0 = 0;
    assign const_716_0 = 0;
    assign const_717_57896044618658097711785492504343953926634992332820282019728792003956564819967 = 57896044618658097711785492504343953926634992332820282019728792003956564819967;
    assign const_719_0 = 0;
    assign const_720_0 = 0;
    assign const_721_0 = 0;
    assign const_722_0 = 0;
    assign const_723_0 = 0;
    assign const_724_0 = 0;
    assign const_725_0 = 0;
    assign const_726_0 = 0;
    assign const_727_0 = 0;
    assign const_728_0 = 0;
    assign const_729_0 = 0;
    assign const_730_0 = 0;
    assign const_731_0 = 0;
    assign const_732_0 = 0;
    assign const_733_0 = 0;
    assign const_734_0 = 0;
    assign const_735_0 = 0;
    assign const_736_0 = 0;
    assign const_737_0 = 0;
    assign const_738_0 = 0;
    assign const_739_0 = 0;
    assign const_740_0 = 0;
    assign const_741_0 = 0;
    assign const_742_0 = 0;
    assign const_743_0 = 0;
    assign const_744_1 = 1;
    assign const_745_0 = 0;
    assign const_746_2 = 2;
    assign const_747_0 = 0;
    assign const_748_3 = 3;
    assign const_749_0 = 0;
    assign const_750_15 = 15;
    assign const_751_0 = 0;
    assign const_752_4 = 4;
    assign const_753_5 = 5;
    assign const_754_6 = 6;
    assign const_755_7 = 7;
    assign const_756_15 = 15;
    assign const_757_0 = 0;
    assign const_758_8 = 8;
    assign const_759_0 = 0;
    assign const_760_6 = 6;
    assign const_761_7 = 7;
    assign const_762_15 = 15;
    assign const_763_0 = 0;
    assign const_764_0 = 0;
    assign const_765_0 = 0;
    assign const_766_1 = 1;
    assign const_767_1 = 1;
    assign const_768_0 = 0;
    assign const_769_1 = 1;
    assign const_770_2 = 2;
    assign const_771_2 = 2;
    assign const_772_0 = 0;
    assign const_773_1 = 1;
    assign const_774_3 = 3;
    assign const_775_3 = 3;
    assign const_776_0 = 0;
    assign const_777_1 = 1;
    assign const_778_0 = 0;
    assign const_779_0 = 0;
    assign const_780_0 = 0;
    assign const_781_0 = 0;
    assign const_782_0 = 0;
    assign const_783_0 = 0;
    assign blue_o = tmp7725;
    assign cfg_speculative_egest = const_0_1;
    assign green_o = tmp7714;
    assign my_calculator_ctrl = tmp7773;
    assign my_calculator_in_x = tmp7776;
    assign my_calculator_in_y = tmp7779;
    assign my_calculator_out_z = tmp7650;
    assign red_o = tmp7703;
    assign tmp1 = {const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0};
    assign tmp2 = {tmp1, const_1_1};
    assign tmp3 = tmp0 + tmp2;
    assign tmp4 = {tmp3[25], tmp3[24], tmp3[23], tmp3[22], tmp3[21], tmp3[20], tmp3[19], tmp3[18], tmp3[17], tmp3[16], tmp3[15], tmp3[14], tmp3[13], tmp3[12], tmp3[11], tmp3[10], tmp3[9], tmp3[8], tmp3[7], tmp3[6], tmp3[5], tmp3[4], tmp3[3], tmp3[2], tmp3[1], tmp3[0]};
    assign tmp6 = {tmp0[24]};
    assign tmp8 = {tmp0[24]};
    assign tmp9 = tmp5 == tmp8;
    assign tmp10 = ~tmp9;
    assign tmp20 = tmp7651;
    assign tmp21 = tmp7652;
    assign tmp22 = tmp7653;
    assign tmp23 = tmp7654;
    assign tmp24 = tmp7655;
    assign tmp25 = tmp7659;
    assign tmp26 = tmp7663;
    assign tmp27 = tmp7667;
    assign tmp28 = tmp7671;
    assign tmp29 = tmp7675;
    assign tmp30 = tmp7679;
    assign tmp31 = tmp7683;
    assign tmp32 = tmp7687;
    assign tmp33 = {const_4_0, const_4_0};
    assign tmp34 = {tmp33, const_3_0};
    assign tmp35 = my_calculator_ctrl == tmp34;
    assign tmp36 = my_calculator_ctrl == const_5_4;
    assign tmp37 = ~tmp35;
    assign tmp38 = tmp37 & tmp36;
    assign tmp39 = ~tmp35;
    assign tmp40 = tmp39 & tmp36;
    assign tmp41 = ~tmp35;
    assign tmp42 = tmp41 & tmp36;
    assign tmp43 = ~tmp35;
    assign tmp44 = tmp43 & tmp36;
    assign tmp45 = ~tmp35;
    assign tmp46 = tmp45 & tmp36;
    assign tmp47 = ~tmp35;
    assign tmp48 = tmp47 & tmp36;
    assign tmp49 = ~tmp35;
    assign tmp50 = tmp49 & tmp36;
    assign tmp51 = ~tmp35;
    assign tmp52 = tmp51 & tmp36;
    assign tmp53 = ~tmp35;
    assign tmp54 = tmp53 & tmp36;
    assign tmp55 = {const_16_0, const_16_0};
    assign tmp56 = {tmp55, const_15_1};
    assign tmp57 = my_calculator_ctrl == tmp56;
    assign tmp58 = ~tmp35;
    assign tmp59 = ~tmp36;
    assign tmp60 = tmp58 & tmp59;
    assign tmp61 = tmp60 & tmp57;
    assign tmp62 = ~tmp35;
    assign tmp63 = ~tmp36;
    assign tmp64 = tmp62 & tmp63;
    assign tmp65 = tmp64 & tmp57;
    assign tmp66 = {const_19_0, const_19_0, const_19_0};
    assign tmp67 = {tmp66, const_18_0};
    assign tmp68 = my_calculator_in_x == tmp67;
    assign tmp69 = my_calculator_in_x == const_20_15;
    assign tmp70 = ~tmp35;
    assign tmp71 = ~tmp36;
    assign tmp72 = tmp70 & tmp71;
    assign tmp73 = tmp72 & tmp57;
    assign tmp74 = ~tmp68;
    assign tmp75 = tmp73 & tmp74;
    assign tmp76 = tmp75 & tmp69;
    assign tmp77 = ~tmp35;
    assign tmp78 = ~tmp36;
    assign tmp79 = tmp77 & tmp78;
    assign tmp80 = tmp79 & tmp57;
    assign tmp81 = ~tmp68;
    assign tmp82 = tmp80 & tmp81;
    assign tmp83 = tmp82 & tmp69;
    assign tmp84 = ~tmp35;
    assign tmp85 = ~tmp36;
    assign tmp86 = tmp84 & tmp85;
    assign tmp87 = tmp86 & tmp57;
    assign tmp88 = ~tmp68;
    assign tmp89 = tmp87 & tmp88;
    assign tmp90 = tmp89 & tmp69;
    assign tmp91 = ~tmp35;
    assign tmp92 = ~tmp36;
    assign tmp93 = tmp91 & tmp92;
    assign tmp94 = tmp93 & tmp57;
    assign tmp95 = ~tmp68;
    assign tmp96 = tmp94 & tmp95;
    assign tmp97 = tmp96 & tmp69;
    assign tmp98 = {const_22_0, const_22_0, const_22_0};
    assign tmp99 = {tmp98, const_21_1};
    assign tmp100 = my_calculator_in_x == tmp99;
    assign tmp101 = {const_24_0, const_24_0};
    assign tmp102 = {tmp101, const_23_2};
    assign tmp103 = my_calculator_in_x == tmp102;
    assign tmp104 = tmp100 | tmp103;
    assign tmp105 = {const_26_0, const_26_0};
    assign tmp106 = {tmp105, const_25_3};
    assign tmp107 = my_calculator_in_x == tmp106;
    assign tmp108 = tmp104 | tmp107;
    assign tmp109 = {tmp11[254], tmp11[253], tmp11[252], tmp11[251], tmp11[250], tmp11[249], tmp11[248], tmp11[247], tmp11[246], tmp11[245], tmp11[244], tmp11[243], tmp11[242], tmp11[241], tmp11[240], tmp11[239], tmp11[238], tmp11[237], tmp11[236], tmp11[235], tmp11[234], tmp11[233], tmp11[232], tmp11[231], tmp11[230], tmp11[229], tmp11[228], tmp11[227], tmp11[226], tmp11[225], tmp11[224], tmp11[223], tmp11[222], tmp11[221], tmp11[220], tmp11[219], tmp11[218], tmp11[217], tmp11[216], tmp11[215], tmp11[214], tmp11[213], tmp11[212], tmp11[211], tmp11[210], tmp11[209], tmp11[208], tmp11[207], tmp11[206], tmp11[205], tmp11[204], tmp11[203], tmp11[202], tmp11[201], tmp11[200], tmp11[199], tmp11[198], tmp11[197], tmp11[196], tmp11[195], tmp11[194], tmp11[193], tmp11[192], tmp11[191], tmp11[190], tmp11[189], tmp11[188], tmp11[187], tmp11[186], tmp11[185], tmp11[184], tmp11[183], tmp11[182], tmp11[181], tmp11[180], tmp11[179], tmp11[178], tmp11[177], tmp11[176], tmp11[175], tmp11[174], tmp11[173], tmp11[172], tmp11[171], tmp11[170], tmp11[169], tmp11[168], tmp11[167], tmp11[166], tmp11[165], tmp11[164], tmp11[163], tmp11[162], tmp11[161], tmp11[160], tmp11[159], tmp11[158], tmp11[157], tmp11[156], tmp11[155], tmp11[154], tmp11[153], tmp11[152], tmp11[151], tmp11[150], tmp11[149], tmp11[148], tmp11[147], tmp11[146], tmp11[145], tmp11[144], tmp11[143], tmp11[142], tmp11[141], tmp11[140], tmp11[139], tmp11[138], tmp11[137], tmp11[136], tmp11[135], tmp11[134], tmp11[133], tmp11[132], tmp11[131], tmp11[130], tmp11[129], tmp11[128], tmp11[127], tmp11[126], tmp11[125], tmp11[124], tmp11[123], tmp11[122], tmp11[121], tmp11[120], tmp11[119], tmp11[118], tmp11[117], tmp11[116], tmp11[115], tmp11[114], tmp11[113], tmp11[112], tmp11[111], tmp11[110], tmp11[109], tmp11[108], tmp11[107], tmp11[106], tmp11[105], tmp11[104], tmp11[103], tmp11[102], tmp11[101], tmp11[100], tmp11[99], tmp11[98], tmp11[97], tmp11[96], tmp11[95], tmp11[94], tmp11[93], tmp11[92], tmp11[91], tmp11[90], tmp11[89], tmp11[88], tmp11[87], tmp11[86], tmp11[85], tmp11[84], tmp11[83], tmp11[82], tmp11[81], tmp11[80], tmp11[79], tmp11[78], tmp11[77], tmp11[76], tmp11[75], tmp11[74], tmp11[73], tmp11[72], tmp11[71], tmp11[70], tmp11[69], tmp11[68], tmp11[67], tmp11[66], tmp11[65], tmp11[64], tmp11[63], tmp11[62], tmp11[61], tmp11[60], tmp11[59], tmp11[58], tmp11[57], tmp11[56], tmp11[55], tmp11[54], tmp11[53], tmp11[52], tmp11[51], tmp11[50], tmp11[49], tmp11[48], tmp11[47], tmp11[46], tmp11[45], tmp11[44], tmp11[43], tmp11[42], tmp11[41], tmp11[40], tmp11[39], tmp11[38], tmp11[37], tmp11[36], tmp11[35], tmp11[34], tmp11[33], tmp11[32], tmp11[31], tmp11[30], tmp11[29], tmp11[28], tmp11[27], tmp11[26], tmp11[25], tmp11[24], tmp11[23], tmp11[22], tmp11[21], tmp11[20], tmp11[19], tmp11[18], tmp11[17], tmp11[16], tmp11[15], tmp11[14], tmp11[13], tmp11[12], tmp11[11], tmp11[10], tmp11[9], tmp11[8], tmp11[7], tmp11[6], tmp11[5], tmp11[4], tmp11[3], tmp11[2], tmp11[1], tmp11[0]};
    assign tmp110 = {tmp109, const_27_0};
    assign tmp111 = {const_28_0};
    assign tmp112 = {tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111, tmp111};
    assign tmp113 = {tmp112, const_28_0};
    assign tmp114 = {tmp11[255]};
    assign tmp115 = tmp113 - tmp11;
    assign tmp116 = {tmp115[256]};
    assign tmp117 = {tmp113[255]};
    assign tmp118 = ~tmp117;
    assign tmp119 = tmp116 ^ tmp118;
    assign tmp120 = {tmp11[255]};
    assign tmp121 = ~tmp120;
    assign tmp122 = tmp119 ^ tmp121;
    assign tmp123 = {tmp110[255]};
    assign tmp124 = {const_29_0};
    assign tmp125 = {tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124, tmp124};
    assign tmp126 = {tmp125, const_29_0};
    assign tmp127 = tmp110 - tmp126;
    assign tmp128 = {tmp127[256]};
    assign tmp129 = {tmp110[255]};
    assign tmp130 = ~tmp129;
    assign tmp131 = tmp128 ^ tmp130;
    assign tmp132 = {tmp126[255]};
    assign tmp133 = ~tmp132;
    assign tmp134 = tmp131 ^ tmp133;
    assign tmp135 = tmp122 & tmp134;
    assign tmp136 = {tmp11[255]};
    assign tmp137 = {const_30_0};
    assign tmp138 = {tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137, tmp137};
    assign tmp139 = {tmp138, const_30_0};
    assign tmp140 = tmp11 - tmp139;
    assign tmp141 = {tmp140[256]};
    assign tmp142 = {tmp11[255]};
    assign tmp143 = ~tmp142;
    assign tmp144 = tmp141 ^ tmp143;
    assign tmp145 = {tmp139[255]};
    assign tmp146 = ~tmp145;
    assign tmp147 = tmp144 ^ tmp146;
    assign tmp148 = {const_31_0};
    assign tmp149 = {tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148, tmp148};
    assign tmp150 = {tmp149, const_31_0};
    assign tmp151 = {tmp110[255]};
    assign tmp152 = tmp150 - tmp110;
    assign tmp153 = {tmp152[256]};
    assign tmp154 = {tmp150[255]};
    assign tmp155 = ~tmp154;
    assign tmp156 = tmp153 ^ tmp155;
    assign tmp157 = {tmp110[255]};
    assign tmp158 = ~tmp157;
    assign tmp159 = tmp156 ^ tmp158;
    assign tmp160 = tmp150 == tmp110;
    assign tmp161 = tmp159 | tmp160;
    assign tmp162 = tmp147 & tmp161;
    assign tmp163 = tmp135 ? const_32_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp110;
    assign tmp164 = tmp162 ? _ver_out_tmp_15 : tmp163;
    assign tmp165 = ~tmp35;
    assign tmp166 = ~tmp36;
    assign tmp167 = tmp165 & tmp166;
    assign tmp168 = tmp167 & tmp57;
    assign tmp169 = ~tmp68;
    assign tmp170 = tmp168 & tmp169;
    assign tmp171 = ~tmp69;
    assign tmp172 = tmp170 & tmp171;
    assign tmp173 = tmp172 & tmp108;
    assign tmp174 = {tmp12[254], tmp12[253], tmp12[252], tmp12[251], tmp12[250], tmp12[249], tmp12[248], tmp12[247], tmp12[246], tmp12[245], tmp12[244], tmp12[243], tmp12[242], tmp12[241], tmp12[240], tmp12[239], tmp12[238], tmp12[237], tmp12[236], tmp12[235], tmp12[234], tmp12[233], tmp12[232], tmp12[231], tmp12[230], tmp12[229], tmp12[228], tmp12[227], tmp12[226], tmp12[225], tmp12[224], tmp12[223], tmp12[222], tmp12[221], tmp12[220], tmp12[219], tmp12[218], tmp12[217], tmp12[216], tmp12[215], tmp12[214], tmp12[213], tmp12[212], tmp12[211], tmp12[210], tmp12[209], tmp12[208], tmp12[207], tmp12[206], tmp12[205], tmp12[204], tmp12[203], tmp12[202], tmp12[201], tmp12[200], tmp12[199], tmp12[198], tmp12[197], tmp12[196], tmp12[195], tmp12[194], tmp12[193], tmp12[192], tmp12[191], tmp12[190], tmp12[189], tmp12[188], tmp12[187], tmp12[186], tmp12[185], tmp12[184], tmp12[183], tmp12[182], tmp12[181], tmp12[180], tmp12[179], tmp12[178], tmp12[177], tmp12[176], tmp12[175], tmp12[174], tmp12[173], tmp12[172], tmp12[171], tmp12[170], tmp12[169], tmp12[168], tmp12[167], tmp12[166], tmp12[165], tmp12[164], tmp12[163], tmp12[162], tmp12[161], tmp12[160], tmp12[159], tmp12[158], tmp12[157], tmp12[156], tmp12[155], tmp12[154], tmp12[153], tmp12[152], tmp12[151], tmp12[150], tmp12[149], tmp12[148], tmp12[147], tmp12[146], tmp12[145], tmp12[144], tmp12[143], tmp12[142], tmp12[141], tmp12[140], tmp12[139], tmp12[138], tmp12[137], tmp12[136], tmp12[135], tmp12[134], tmp12[133], tmp12[132], tmp12[131], tmp12[130], tmp12[129], tmp12[128], tmp12[127], tmp12[126], tmp12[125], tmp12[124], tmp12[123], tmp12[122], tmp12[121], tmp12[120], tmp12[119], tmp12[118], tmp12[117], tmp12[116], tmp12[115], tmp12[114], tmp12[113], tmp12[112], tmp12[111], tmp12[110], tmp12[109], tmp12[108], tmp12[107], tmp12[106], tmp12[105], tmp12[104], tmp12[103], tmp12[102], tmp12[101], tmp12[100], tmp12[99], tmp12[98], tmp12[97], tmp12[96], tmp12[95], tmp12[94], tmp12[93], tmp12[92], tmp12[91], tmp12[90], tmp12[89], tmp12[88], tmp12[87], tmp12[86], tmp12[85], tmp12[84], tmp12[83], tmp12[82], tmp12[81], tmp12[80], tmp12[79], tmp12[78], tmp12[77], tmp12[76], tmp12[75], tmp12[74], tmp12[73], tmp12[72], tmp12[71], tmp12[70], tmp12[69], tmp12[68], tmp12[67], tmp12[66], tmp12[65], tmp12[64], tmp12[63], tmp12[62], tmp12[61], tmp12[60], tmp12[59], tmp12[58], tmp12[57], tmp12[56], tmp12[55], tmp12[54], tmp12[53], tmp12[52], tmp12[51], tmp12[50], tmp12[49], tmp12[48], tmp12[47], tmp12[46], tmp12[45], tmp12[44], tmp12[43], tmp12[42], tmp12[41], tmp12[40], tmp12[39], tmp12[38], tmp12[37], tmp12[36], tmp12[35], tmp12[34], tmp12[33], tmp12[32], tmp12[31], tmp12[30], tmp12[29], tmp12[28], tmp12[27], tmp12[26], tmp12[25], tmp12[24], tmp12[23], tmp12[22], tmp12[21], tmp12[20], tmp12[19], tmp12[18], tmp12[17], tmp12[16], tmp12[15], tmp12[14], tmp12[13], tmp12[12], tmp12[11], tmp12[10], tmp12[9], tmp12[8], tmp12[7], tmp12[6], tmp12[5], tmp12[4], tmp12[3], tmp12[2], tmp12[1], tmp12[0]};
    assign tmp175 = {tmp174, const_34_0};
    assign tmp176 = {const_35_0};
    assign tmp177 = {tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176, tmp176};
    assign tmp178 = {tmp177, const_35_0};
    assign tmp179 = {tmp12[255]};
    assign tmp180 = tmp178 - tmp12;
    assign tmp181 = {tmp180[256]};
    assign tmp182 = {tmp178[255]};
    assign tmp183 = ~tmp182;
    assign tmp184 = tmp181 ^ tmp183;
    assign tmp185 = {tmp12[255]};
    assign tmp186 = ~tmp185;
    assign tmp187 = tmp184 ^ tmp186;
    assign tmp188 = {tmp175[255]};
    assign tmp189 = {const_36_0};
    assign tmp190 = {tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189, tmp189};
    assign tmp191 = {tmp190, const_36_0};
    assign tmp192 = tmp175 - tmp191;
    assign tmp193 = {tmp192[256]};
    assign tmp194 = {tmp175[255]};
    assign tmp195 = ~tmp194;
    assign tmp196 = tmp193 ^ tmp195;
    assign tmp197 = {tmp191[255]};
    assign tmp198 = ~tmp197;
    assign tmp199 = tmp196 ^ tmp198;
    assign tmp200 = tmp187 & tmp199;
    assign tmp201 = {tmp12[255]};
    assign tmp202 = {const_37_0};
    assign tmp203 = {tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202, tmp202};
    assign tmp204 = {tmp203, const_37_0};
    assign tmp205 = tmp12 - tmp204;
    assign tmp206 = {tmp205[256]};
    assign tmp207 = {tmp12[255]};
    assign tmp208 = ~tmp207;
    assign tmp209 = tmp206 ^ tmp208;
    assign tmp210 = {tmp204[255]};
    assign tmp211 = ~tmp210;
    assign tmp212 = tmp209 ^ tmp211;
    assign tmp213 = {const_38_0};
    assign tmp214 = {tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213, tmp213};
    assign tmp215 = {tmp214, const_38_0};
    assign tmp216 = {tmp175[255]};
    assign tmp217 = tmp215 - tmp175;
    assign tmp218 = {tmp217[256]};
    assign tmp219 = {tmp215[255]};
    assign tmp220 = ~tmp219;
    assign tmp221 = tmp218 ^ tmp220;
    assign tmp222 = {tmp175[255]};
    assign tmp223 = ~tmp222;
    assign tmp224 = tmp221 ^ tmp223;
    assign tmp225 = tmp215 == tmp175;
    assign tmp226 = tmp224 | tmp225;
    assign tmp227 = tmp212 & tmp226;
    assign tmp228 = tmp200 ? const_39_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp175;
    assign tmp229 = tmp227 ? _ver_out_tmp_19 : tmp228;
    assign tmp230 = ~tmp35;
    assign tmp231 = ~tmp36;
    assign tmp232 = tmp230 & tmp231;
    assign tmp233 = tmp232 & tmp57;
    assign tmp234 = ~tmp68;
    assign tmp235 = tmp233 & tmp234;
    assign tmp236 = ~tmp69;
    assign tmp237 = tmp235 & tmp236;
    assign tmp238 = tmp237 & tmp108;
    assign tmp239 = {tmp15[254], tmp15[253], tmp15[252], tmp15[251], tmp15[250], tmp15[249], tmp15[248], tmp15[247], tmp15[246], tmp15[245], tmp15[244], tmp15[243], tmp15[242], tmp15[241], tmp15[240], tmp15[239], tmp15[238], tmp15[237], tmp15[236], tmp15[235], tmp15[234], tmp15[233], tmp15[232], tmp15[231], tmp15[230], tmp15[229], tmp15[228], tmp15[227], tmp15[226], tmp15[225], tmp15[224], tmp15[223], tmp15[222], tmp15[221], tmp15[220], tmp15[219], tmp15[218], tmp15[217], tmp15[216], tmp15[215], tmp15[214], tmp15[213], tmp15[212], tmp15[211], tmp15[210], tmp15[209], tmp15[208], tmp15[207], tmp15[206], tmp15[205], tmp15[204], tmp15[203], tmp15[202], tmp15[201], tmp15[200], tmp15[199], tmp15[198], tmp15[197], tmp15[196], tmp15[195], tmp15[194], tmp15[193], tmp15[192], tmp15[191], tmp15[190], tmp15[189], tmp15[188], tmp15[187], tmp15[186], tmp15[185], tmp15[184], tmp15[183], tmp15[182], tmp15[181], tmp15[180], tmp15[179], tmp15[178], tmp15[177], tmp15[176], tmp15[175], tmp15[174], tmp15[173], tmp15[172], tmp15[171], tmp15[170], tmp15[169], tmp15[168], tmp15[167], tmp15[166], tmp15[165], tmp15[164], tmp15[163], tmp15[162], tmp15[161], tmp15[160], tmp15[159], tmp15[158], tmp15[157], tmp15[156], tmp15[155], tmp15[154], tmp15[153], tmp15[152], tmp15[151], tmp15[150], tmp15[149], tmp15[148], tmp15[147], tmp15[146], tmp15[145], tmp15[144], tmp15[143], tmp15[142], tmp15[141], tmp15[140], tmp15[139], tmp15[138], tmp15[137], tmp15[136], tmp15[135], tmp15[134], tmp15[133], tmp15[132], tmp15[131], tmp15[130], tmp15[129], tmp15[128], tmp15[127], tmp15[126], tmp15[125], tmp15[124], tmp15[123], tmp15[122], tmp15[121], tmp15[120], tmp15[119], tmp15[118], tmp15[117], tmp15[116], tmp15[115], tmp15[114], tmp15[113], tmp15[112], tmp15[111], tmp15[110], tmp15[109], tmp15[108], tmp15[107], tmp15[106], tmp15[105], tmp15[104], tmp15[103], tmp15[102], tmp15[101], tmp15[100], tmp15[99], tmp15[98], tmp15[97], tmp15[96], tmp15[95], tmp15[94], tmp15[93], tmp15[92], tmp15[91], tmp15[90], tmp15[89], tmp15[88], tmp15[87], tmp15[86], tmp15[85], tmp15[84], tmp15[83], tmp15[82], tmp15[81], tmp15[80], tmp15[79], tmp15[78], tmp15[77], tmp15[76], tmp15[75], tmp15[74], tmp15[73], tmp15[72], tmp15[71], tmp15[70], tmp15[69], tmp15[68], tmp15[67], tmp15[66], tmp15[65], tmp15[64], tmp15[63], tmp15[62], tmp15[61], tmp15[60], tmp15[59], tmp15[58], tmp15[57], tmp15[56], tmp15[55], tmp15[54], tmp15[53], tmp15[52], tmp15[51], tmp15[50], tmp15[49], tmp15[48], tmp15[47], tmp15[46], tmp15[45], tmp15[44], tmp15[43], tmp15[42], tmp15[41], tmp15[40], tmp15[39], tmp15[38], tmp15[37], tmp15[36], tmp15[35], tmp15[34], tmp15[33], tmp15[32], tmp15[31], tmp15[30], tmp15[29], tmp15[28], tmp15[27], tmp15[26], tmp15[25], tmp15[24], tmp15[23], tmp15[22], tmp15[21], tmp15[20], tmp15[19], tmp15[18], tmp15[17], tmp15[16], tmp15[15], tmp15[14], tmp15[13], tmp15[12], tmp15[11], tmp15[10], tmp15[9], tmp15[8], tmp15[7], tmp15[6], tmp15[5], tmp15[4], tmp15[3], tmp15[2], tmp15[1], tmp15[0]};
    assign tmp240 = {tmp239, const_41_0};
    assign tmp241 = {const_42_0};
    assign tmp242 = {tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241, tmp241};
    assign tmp243 = {tmp242, const_42_0};
    assign tmp244 = {tmp15[255]};
    assign tmp245 = tmp243 - tmp15;
    assign tmp246 = {tmp245[256]};
    assign tmp247 = {tmp243[255]};
    assign tmp248 = ~tmp247;
    assign tmp249 = tmp246 ^ tmp248;
    assign tmp250 = {tmp15[255]};
    assign tmp251 = ~tmp250;
    assign tmp252 = tmp249 ^ tmp251;
    assign tmp253 = {tmp240[255]};
    assign tmp254 = {const_43_0};
    assign tmp255 = {tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254, tmp254};
    assign tmp256 = {tmp255, const_43_0};
    assign tmp257 = tmp240 - tmp256;
    assign tmp258 = {tmp257[256]};
    assign tmp259 = {tmp240[255]};
    assign tmp260 = ~tmp259;
    assign tmp261 = tmp258 ^ tmp260;
    assign tmp262 = {tmp256[255]};
    assign tmp263 = ~tmp262;
    assign tmp264 = tmp261 ^ tmp263;
    assign tmp265 = tmp252 & tmp264;
    assign tmp266 = {tmp15[255]};
    assign tmp267 = {const_44_0};
    assign tmp268 = {tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267, tmp267};
    assign tmp269 = {tmp268, const_44_0};
    assign tmp270 = tmp15 - tmp269;
    assign tmp271 = {tmp270[256]};
    assign tmp272 = {tmp15[255]};
    assign tmp273 = ~tmp272;
    assign tmp274 = tmp271 ^ tmp273;
    assign tmp275 = {tmp269[255]};
    assign tmp276 = ~tmp275;
    assign tmp277 = tmp274 ^ tmp276;
    assign tmp278 = {const_45_0};
    assign tmp279 = {tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278, tmp278};
    assign tmp280 = {tmp279, const_45_0};
    assign tmp281 = {tmp240[255]};
    assign tmp282 = tmp280 - tmp240;
    assign tmp283 = {tmp282[256]};
    assign tmp284 = {tmp280[255]};
    assign tmp285 = ~tmp284;
    assign tmp286 = tmp283 ^ tmp285;
    assign tmp287 = {tmp240[255]};
    assign tmp288 = ~tmp287;
    assign tmp289 = tmp286 ^ tmp288;
    assign tmp290 = tmp280 == tmp240;
    assign tmp291 = tmp289 | tmp290;
    assign tmp292 = tmp277 & tmp291;
    assign tmp293 = tmp265 ? const_46_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp240;
    assign tmp294 = tmp292 ? _ver_out_tmp_22 : tmp293;
    assign tmp295 = ~tmp35;
    assign tmp296 = ~tmp36;
    assign tmp297 = tmp295 & tmp296;
    assign tmp298 = tmp297 & tmp57;
    assign tmp299 = ~tmp68;
    assign tmp300 = tmp298 & tmp299;
    assign tmp301 = ~tmp69;
    assign tmp302 = tmp300 & tmp301;
    assign tmp303 = tmp302 & tmp108;
    assign tmp304 = {tmp16[254], tmp16[253], tmp16[252], tmp16[251], tmp16[250], tmp16[249], tmp16[248], tmp16[247], tmp16[246], tmp16[245], tmp16[244], tmp16[243], tmp16[242], tmp16[241], tmp16[240], tmp16[239], tmp16[238], tmp16[237], tmp16[236], tmp16[235], tmp16[234], tmp16[233], tmp16[232], tmp16[231], tmp16[230], tmp16[229], tmp16[228], tmp16[227], tmp16[226], tmp16[225], tmp16[224], tmp16[223], tmp16[222], tmp16[221], tmp16[220], tmp16[219], tmp16[218], tmp16[217], tmp16[216], tmp16[215], tmp16[214], tmp16[213], tmp16[212], tmp16[211], tmp16[210], tmp16[209], tmp16[208], tmp16[207], tmp16[206], tmp16[205], tmp16[204], tmp16[203], tmp16[202], tmp16[201], tmp16[200], tmp16[199], tmp16[198], tmp16[197], tmp16[196], tmp16[195], tmp16[194], tmp16[193], tmp16[192], tmp16[191], tmp16[190], tmp16[189], tmp16[188], tmp16[187], tmp16[186], tmp16[185], tmp16[184], tmp16[183], tmp16[182], tmp16[181], tmp16[180], tmp16[179], tmp16[178], tmp16[177], tmp16[176], tmp16[175], tmp16[174], tmp16[173], tmp16[172], tmp16[171], tmp16[170], tmp16[169], tmp16[168], tmp16[167], tmp16[166], tmp16[165], tmp16[164], tmp16[163], tmp16[162], tmp16[161], tmp16[160], tmp16[159], tmp16[158], tmp16[157], tmp16[156], tmp16[155], tmp16[154], tmp16[153], tmp16[152], tmp16[151], tmp16[150], tmp16[149], tmp16[148], tmp16[147], tmp16[146], tmp16[145], tmp16[144], tmp16[143], tmp16[142], tmp16[141], tmp16[140], tmp16[139], tmp16[138], tmp16[137], tmp16[136], tmp16[135], tmp16[134], tmp16[133], tmp16[132], tmp16[131], tmp16[130], tmp16[129], tmp16[128], tmp16[127], tmp16[126], tmp16[125], tmp16[124], tmp16[123], tmp16[122], tmp16[121], tmp16[120], tmp16[119], tmp16[118], tmp16[117], tmp16[116], tmp16[115], tmp16[114], tmp16[113], tmp16[112], tmp16[111], tmp16[110], tmp16[109], tmp16[108], tmp16[107], tmp16[106], tmp16[105], tmp16[104], tmp16[103], tmp16[102], tmp16[101], tmp16[100], tmp16[99], tmp16[98], tmp16[97], tmp16[96], tmp16[95], tmp16[94], tmp16[93], tmp16[92], tmp16[91], tmp16[90], tmp16[89], tmp16[88], tmp16[87], tmp16[86], tmp16[85], tmp16[84], tmp16[83], tmp16[82], tmp16[81], tmp16[80], tmp16[79], tmp16[78], tmp16[77], tmp16[76], tmp16[75], tmp16[74], tmp16[73], tmp16[72], tmp16[71], tmp16[70], tmp16[69], tmp16[68], tmp16[67], tmp16[66], tmp16[65], tmp16[64], tmp16[63], tmp16[62], tmp16[61], tmp16[60], tmp16[59], tmp16[58], tmp16[57], tmp16[56], tmp16[55], tmp16[54], tmp16[53], tmp16[52], tmp16[51], tmp16[50], tmp16[49], tmp16[48], tmp16[47], tmp16[46], tmp16[45], tmp16[44], tmp16[43], tmp16[42], tmp16[41], tmp16[40], tmp16[39], tmp16[38], tmp16[37], tmp16[36], tmp16[35], tmp16[34], tmp16[33], tmp16[32], tmp16[31], tmp16[30], tmp16[29], tmp16[28], tmp16[27], tmp16[26], tmp16[25], tmp16[24], tmp16[23], tmp16[22], tmp16[21], tmp16[20], tmp16[19], tmp16[18], tmp16[17], tmp16[16], tmp16[15], tmp16[14], tmp16[13], tmp16[12], tmp16[11], tmp16[10], tmp16[9], tmp16[8], tmp16[7], tmp16[6], tmp16[5], tmp16[4], tmp16[3], tmp16[2], tmp16[1], tmp16[0]};
    assign tmp305 = {tmp304, const_48_0};
    assign tmp306 = {const_49_0};
    assign tmp307 = {tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306, tmp306};
    assign tmp308 = {tmp307, const_49_0};
    assign tmp309 = {tmp16[255]};
    assign tmp310 = tmp308 - tmp16;
    assign tmp311 = {tmp310[256]};
    assign tmp312 = {tmp308[255]};
    assign tmp313 = ~tmp312;
    assign tmp314 = tmp311 ^ tmp313;
    assign tmp315 = {tmp16[255]};
    assign tmp316 = ~tmp315;
    assign tmp317 = tmp314 ^ tmp316;
    assign tmp318 = {tmp305[255]};
    assign tmp319 = {const_50_0};
    assign tmp320 = {tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319, tmp319};
    assign tmp321 = {tmp320, const_50_0};
    assign tmp322 = tmp305 - tmp321;
    assign tmp323 = {tmp322[256]};
    assign tmp324 = {tmp305[255]};
    assign tmp325 = ~tmp324;
    assign tmp326 = tmp323 ^ tmp325;
    assign tmp327 = {tmp321[255]};
    assign tmp328 = ~tmp327;
    assign tmp329 = tmp326 ^ tmp328;
    assign tmp330 = tmp317 & tmp329;
    assign tmp331 = {tmp16[255]};
    assign tmp332 = {const_51_0};
    assign tmp333 = {tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332, tmp332};
    assign tmp334 = {tmp333, const_51_0};
    assign tmp335 = tmp16 - tmp334;
    assign tmp336 = {tmp335[256]};
    assign tmp337 = {tmp16[255]};
    assign tmp338 = ~tmp337;
    assign tmp339 = tmp336 ^ tmp338;
    assign tmp340 = {tmp334[255]};
    assign tmp341 = ~tmp340;
    assign tmp342 = tmp339 ^ tmp341;
    assign tmp343 = {const_52_0};
    assign tmp344 = {tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343, tmp343};
    assign tmp345 = {tmp344, const_52_0};
    assign tmp346 = {tmp305[255]};
    assign tmp347 = tmp345 - tmp305;
    assign tmp348 = {tmp347[256]};
    assign tmp349 = {tmp345[255]};
    assign tmp350 = ~tmp349;
    assign tmp351 = tmp348 ^ tmp350;
    assign tmp352 = {tmp305[255]};
    assign tmp353 = ~tmp352;
    assign tmp354 = tmp351 ^ tmp353;
    assign tmp355 = tmp345 == tmp305;
    assign tmp356 = tmp354 | tmp355;
    assign tmp357 = tmp342 & tmp356;
    assign tmp358 = tmp330 ? const_53_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp305;
    assign tmp359 = tmp357 ? _ver_out_tmp_24 : tmp358;
    assign tmp360 = ~tmp35;
    assign tmp361 = ~tmp36;
    assign tmp362 = tmp360 & tmp361;
    assign tmp363 = tmp362 & tmp57;
    assign tmp364 = ~tmp68;
    assign tmp365 = tmp363 & tmp364;
    assign tmp366 = ~tmp69;
    assign tmp367 = tmp365 & tmp366;
    assign tmp368 = tmp367 & tmp108;
    assign tmp369 = {const_56_0};
    assign tmp370 = {tmp369, const_55_6};
    assign tmp371 = my_calculator_in_x == tmp370;
    assign tmp372 = {const_58_0};
    assign tmp373 = {tmp372, const_57_7};
    assign tmp374 = my_calculator_in_x == tmp373;
    assign tmp375 = tmp371 | tmp374;
    assign tmp376 = ~tmp35;
    assign tmp377 = ~tmp36;
    assign tmp378 = tmp376 & tmp377;
    assign tmp379 = tmp378 & tmp57;
    assign tmp380 = ~tmp68;
    assign tmp381 = tmp379 & tmp380;
    assign tmp382 = ~tmp69;
    assign tmp383 = tmp381 & tmp382;
    assign tmp384 = ~tmp108;
    assign tmp385 = tmp383 & tmp384;
    assign tmp386 = tmp385 & tmp375;
    assign tmp387 = ~tmp35;
    assign tmp388 = ~tmp36;
    assign tmp389 = tmp387 & tmp388;
    assign tmp390 = tmp389 & tmp57;
    assign tmp391 = ~tmp68;
    assign tmp392 = tmp390 & tmp391;
    assign tmp393 = ~tmp69;
    assign tmp394 = tmp392 & tmp393;
    assign tmp395 = ~tmp108;
    assign tmp396 = tmp394 & tmp395;
    assign tmp397 = tmp396 & tmp375;
    assign tmp398 = ~tmp35;
    assign tmp399 = ~tmp36;
    assign tmp400 = tmp398 & tmp399;
    assign tmp401 = tmp400 & tmp57;
    assign tmp402 = ~tmp68;
    assign tmp403 = tmp401 & tmp402;
    assign tmp404 = ~tmp69;
    assign tmp405 = tmp403 & tmp404;
    assign tmp406 = ~tmp108;
    assign tmp407 = tmp405 & tmp406;
    assign tmp408 = tmp407 & tmp375;
    assign tmp409 = ~tmp35;
    assign tmp410 = ~tmp36;
    assign tmp411 = tmp409 & tmp410;
    assign tmp412 = tmp411 & tmp57;
    assign tmp413 = ~tmp68;
    assign tmp414 = tmp412 & tmp413;
    assign tmp415 = ~tmp69;
    assign tmp416 = tmp414 & tmp415;
    assign tmp417 = ~tmp108;
    assign tmp418 = tmp416 & tmp417;
    assign tmp419 = tmp418 & tmp375;
    assign tmp420 = ~tmp35;
    assign tmp421 = ~tmp36;
    assign tmp422 = tmp420 & tmp421;
    assign tmp423 = tmp422 & tmp57;
    assign tmp424 = ~tmp68;
    assign tmp425 = tmp423 & tmp424;
    assign tmp426 = ~tmp69;
    assign tmp427 = tmp425 & tmp426;
    assign tmp428 = ~tmp108;
    assign tmp429 = tmp427 & tmp428;
    assign tmp430 = tmp429 & tmp375;
    assign tmp431 = ~tmp35;
    assign tmp432 = ~tmp36;
    assign tmp433 = tmp431 & tmp432;
    assign tmp434 = tmp433 & tmp57;
    assign tmp435 = ~tmp68;
    assign tmp436 = tmp434 & tmp435;
    assign tmp437 = ~tmp69;
    assign tmp438 = tmp436 & tmp437;
    assign tmp439 = ~tmp108;
    assign tmp440 = tmp438 & tmp439;
    assign tmp441 = tmp440 & tmp375;
    assign tmp442 = ~tmp35;
    assign tmp443 = ~tmp36;
    assign tmp444 = tmp442 & tmp443;
    assign tmp445 = tmp444 & tmp57;
    assign tmp446 = ~tmp68;
    assign tmp447 = tmp445 & tmp446;
    assign tmp448 = ~tmp69;
    assign tmp449 = tmp447 & tmp448;
    assign tmp450 = ~tmp108;
    assign tmp451 = tmp449 & tmp450;
    assign tmp452 = tmp451 & tmp375;
    assign tmp453 = ~tmp35;
    assign tmp454 = ~tmp36;
    assign tmp455 = tmp453 & tmp454;
    assign tmp456 = tmp455 & tmp57;
    assign tmp457 = ~tmp68;
    assign tmp458 = tmp456 & tmp457;
    assign tmp459 = ~tmp69;
    assign tmp460 = tmp458 & tmp459;
    assign tmp461 = ~tmp108;
    assign tmp462 = tmp460 & tmp461;
    assign tmp463 = tmp462 & tmp375;
    assign tmp464 = {const_60_0};
    assign tmp465 = {tmp464, const_59_4};
    assign tmp466 = my_calculator_in_x == tmp465;
    assign tmp467 = {const_62_0};
    assign tmp468 = {tmp467, const_61_5};
    assign tmp469 = my_calculator_in_x == tmp468;
    assign tmp470 = tmp466 | tmp469;
    assign tmp471 = {tmp11[255]};
    assign tmp472 = {tmp471};
    assign tmp473 = {tmp472, tmp11};
    assign tmp474 = {tmp13[255]};
    assign tmp475 = {tmp474};
    assign tmp476 = {tmp475, tmp13};
    assign tmp477 = tmp473 + tmp476;
    assign tmp478 = {tmp477[256], tmp477[255], tmp477[254], tmp477[253], tmp477[252], tmp477[251], tmp477[250], tmp477[249], tmp477[248], tmp477[247], tmp477[246], tmp477[245], tmp477[244], tmp477[243], tmp477[242], tmp477[241], tmp477[240], tmp477[239], tmp477[238], tmp477[237], tmp477[236], tmp477[235], tmp477[234], tmp477[233], tmp477[232], tmp477[231], tmp477[230], tmp477[229], tmp477[228], tmp477[227], tmp477[226], tmp477[225], tmp477[224], tmp477[223], tmp477[222], tmp477[221], tmp477[220], tmp477[219], tmp477[218], tmp477[217], tmp477[216], tmp477[215], tmp477[214], tmp477[213], tmp477[212], tmp477[211], tmp477[210], tmp477[209], tmp477[208], tmp477[207], tmp477[206], tmp477[205], tmp477[204], tmp477[203], tmp477[202], tmp477[201], tmp477[200], tmp477[199], tmp477[198], tmp477[197], tmp477[196], tmp477[195], tmp477[194], tmp477[193], tmp477[192], tmp477[191], tmp477[190], tmp477[189], tmp477[188], tmp477[187], tmp477[186], tmp477[185], tmp477[184], tmp477[183], tmp477[182], tmp477[181], tmp477[180], tmp477[179], tmp477[178], tmp477[177], tmp477[176], tmp477[175], tmp477[174], tmp477[173], tmp477[172], tmp477[171], tmp477[170], tmp477[169], tmp477[168], tmp477[167], tmp477[166], tmp477[165], tmp477[164], tmp477[163], tmp477[162], tmp477[161], tmp477[160], tmp477[159], tmp477[158], tmp477[157], tmp477[156], tmp477[155], tmp477[154], tmp477[153], tmp477[152], tmp477[151], tmp477[150], tmp477[149], tmp477[148], tmp477[147], tmp477[146], tmp477[145], tmp477[144], tmp477[143], tmp477[142], tmp477[141], tmp477[140], tmp477[139], tmp477[138], tmp477[137], tmp477[136], tmp477[135], tmp477[134], tmp477[133], tmp477[132], tmp477[131], tmp477[130], tmp477[129], tmp477[128], tmp477[127], tmp477[126], tmp477[125], tmp477[124], tmp477[123], tmp477[122], tmp477[121], tmp477[120], tmp477[119], tmp477[118], tmp477[117], tmp477[116], tmp477[115], tmp477[114], tmp477[113], tmp477[112], tmp477[111], tmp477[110], tmp477[109], tmp477[108], tmp477[107], tmp477[106], tmp477[105], tmp477[104], tmp477[103], tmp477[102], tmp477[101], tmp477[100], tmp477[99], tmp477[98], tmp477[97], tmp477[96], tmp477[95], tmp477[94], tmp477[93], tmp477[92], tmp477[91], tmp477[90], tmp477[89], tmp477[88], tmp477[87], tmp477[86], tmp477[85], tmp477[84], tmp477[83], tmp477[82], tmp477[81], tmp477[80], tmp477[79], tmp477[78], tmp477[77], tmp477[76], tmp477[75], tmp477[74], tmp477[73], tmp477[72], tmp477[71], tmp477[70], tmp477[69], tmp477[68], tmp477[67], tmp477[66], tmp477[65], tmp477[64], tmp477[63], tmp477[62], tmp477[61], tmp477[60], tmp477[59], tmp477[58], tmp477[57], tmp477[56], tmp477[55], tmp477[54], tmp477[53], tmp477[52], tmp477[51], tmp477[50], tmp477[49], tmp477[48], tmp477[47], tmp477[46], tmp477[45], tmp477[44], tmp477[43], tmp477[42], tmp477[41], tmp477[40], tmp477[39], tmp477[38], tmp477[37], tmp477[36], tmp477[35], tmp477[34], tmp477[33], tmp477[32], tmp477[31], tmp477[30], tmp477[29], tmp477[28], tmp477[27], tmp477[26], tmp477[25], tmp477[24], tmp477[23], tmp477[22], tmp477[21], tmp477[20], tmp477[19], tmp477[18], tmp477[17], tmp477[16], tmp477[15], tmp477[14], tmp477[13], tmp477[12], tmp477[11], tmp477[10], tmp477[9], tmp477[8], tmp477[7], tmp477[6], tmp477[5], tmp477[4], tmp477[3], tmp477[2], tmp477[1], tmp477[0]};
    assign tmp479 = {tmp478[255], tmp478[254], tmp478[253], tmp478[252], tmp478[251], tmp478[250], tmp478[249], tmp478[248], tmp478[247], tmp478[246], tmp478[245], tmp478[244], tmp478[243], tmp478[242], tmp478[241], tmp478[240], tmp478[239], tmp478[238], tmp478[237], tmp478[236], tmp478[235], tmp478[234], tmp478[233], tmp478[232], tmp478[231], tmp478[230], tmp478[229], tmp478[228], tmp478[227], tmp478[226], tmp478[225], tmp478[224], tmp478[223], tmp478[222], tmp478[221], tmp478[220], tmp478[219], tmp478[218], tmp478[217], tmp478[216], tmp478[215], tmp478[214], tmp478[213], tmp478[212], tmp478[211], tmp478[210], tmp478[209], tmp478[208], tmp478[207], tmp478[206], tmp478[205], tmp478[204], tmp478[203], tmp478[202], tmp478[201], tmp478[200], tmp478[199], tmp478[198], tmp478[197], tmp478[196], tmp478[195], tmp478[194], tmp478[193], tmp478[192], tmp478[191], tmp478[190], tmp478[189], tmp478[188], tmp478[187], tmp478[186], tmp478[185], tmp478[184], tmp478[183], tmp478[182], tmp478[181], tmp478[180], tmp478[179], tmp478[178], tmp478[177], tmp478[176], tmp478[175], tmp478[174], tmp478[173], tmp478[172], tmp478[171], tmp478[170], tmp478[169], tmp478[168], tmp478[167], tmp478[166], tmp478[165], tmp478[164], tmp478[163], tmp478[162], tmp478[161], tmp478[160], tmp478[159], tmp478[158], tmp478[157], tmp478[156], tmp478[155], tmp478[154], tmp478[153], tmp478[152], tmp478[151], tmp478[150], tmp478[149], tmp478[148], tmp478[147], tmp478[146], tmp478[145], tmp478[144], tmp478[143], tmp478[142], tmp478[141], tmp478[140], tmp478[139], tmp478[138], tmp478[137], tmp478[136], tmp478[135], tmp478[134], tmp478[133], tmp478[132], tmp478[131], tmp478[130], tmp478[129], tmp478[128], tmp478[127], tmp478[126], tmp478[125], tmp478[124], tmp478[123], tmp478[122], tmp478[121], tmp478[120], tmp478[119], tmp478[118], tmp478[117], tmp478[116], tmp478[115], tmp478[114], tmp478[113], tmp478[112], tmp478[111], tmp478[110], tmp478[109], tmp478[108], tmp478[107], tmp478[106], tmp478[105], tmp478[104], tmp478[103], tmp478[102], tmp478[101], tmp478[100], tmp478[99], tmp478[98], tmp478[97], tmp478[96], tmp478[95], tmp478[94], tmp478[93], tmp478[92], tmp478[91], tmp478[90], tmp478[89], tmp478[88], tmp478[87], tmp478[86], tmp478[85], tmp478[84], tmp478[83], tmp478[82], tmp478[81], tmp478[80], tmp478[79], tmp478[78], tmp478[77], tmp478[76], tmp478[75], tmp478[74], tmp478[73], tmp478[72], tmp478[71], tmp478[70], tmp478[69], tmp478[68], tmp478[67], tmp478[66], tmp478[65], tmp478[64], tmp478[63], tmp478[62], tmp478[61], tmp478[60], tmp478[59], tmp478[58], tmp478[57], tmp478[56], tmp478[55], tmp478[54], tmp478[53], tmp478[52], tmp478[51], tmp478[50], tmp478[49], tmp478[48], tmp478[47], tmp478[46], tmp478[45], tmp478[44], tmp478[43], tmp478[42], tmp478[41], tmp478[40], tmp478[39], tmp478[38], tmp478[37], tmp478[36], tmp478[35], tmp478[34], tmp478[33], tmp478[32], tmp478[31], tmp478[30], tmp478[29], tmp478[28], tmp478[27], tmp478[26], tmp478[25], tmp478[24], tmp478[23], tmp478[22], tmp478[21], tmp478[20], tmp478[19], tmp478[18], tmp478[17], tmp478[16], tmp478[15], tmp478[14], tmp478[13], tmp478[12], tmp478[11], tmp478[10], tmp478[9], tmp478[8], tmp478[7], tmp478[6], tmp478[5], tmp478[4], tmp478[3], tmp478[2], tmp478[1], tmp478[0]};
    assign tmp480 = {const_63_0};
    assign tmp481 = {tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480, tmp480};
    assign tmp482 = {tmp481, const_63_0};
    assign tmp483 = {tmp11[255]};
    assign tmp484 = tmp482 - tmp11;
    assign tmp485 = {tmp484[256]};
    assign tmp486 = {tmp482[255]};
    assign tmp487 = ~tmp486;
    assign tmp488 = tmp485 ^ tmp487;
    assign tmp489 = {tmp11[255]};
    assign tmp490 = ~tmp489;
    assign tmp491 = tmp488 ^ tmp490;
    assign tmp492 = {const_64_0};
    assign tmp493 = {tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492, tmp492};
    assign tmp494 = {tmp493, const_64_0};
    assign tmp495 = {tmp13[255]};
    assign tmp496 = tmp494 - tmp13;
    assign tmp497 = {tmp496[256]};
    assign tmp498 = {tmp494[255]};
    assign tmp499 = ~tmp498;
    assign tmp500 = tmp497 ^ tmp499;
    assign tmp501 = {tmp13[255]};
    assign tmp502 = ~tmp501;
    assign tmp503 = tmp500 ^ tmp502;
    assign tmp504 = tmp491 & tmp503;
    assign tmp505 = {tmp479[255]};
    assign tmp506 = {const_65_0};
    assign tmp507 = {tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506, tmp506};
    assign tmp508 = {tmp507, const_65_0};
    assign tmp509 = tmp479 - tmp508;
    assign tmp510 = {tmp509[256]};
    assign tmp511 = {tmp479[255]};
    assign tmp512 = ~tmp511;
    assign tmp513 = tmp510 ^ tmp512;
    assign tmp514 = {tmp508[255]};
    assign tmp515 = ~tmp514;
    assign tmp516 = tmp513 ^ tmp515;
    assign tmp517 = tmp479 == tmp508;
    assign tmp518 = tmp516 | tmp517;
    assign tmp519 = tmp504 & tmp518;
    assign tmp520 = {tmp11[255]};
    assign tmp521 = {const_66_0};
    assign tmp522 = {tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521, tmp521};
    assign tmp523 = {tmp522, const_66_0};
    assign tmp524 = tmp11 - tmp523;
    assign tmp525 = {tmp524[256]};
    assign tmp526 = {tmp11[255]};
    assign tmp527 = ~tmp526;
    assign tmp528 = tmp525 ^ tmp527;
    assign tmp529 = {tmp523[255]};
    assign tmp530 = ~tmp529;
    assign tmp531 = tmp528 ^ tmp530;
    assign tmp532 = {tmp13[255]};
    assign tmp533 = {const_67_0};
    assign tmp534 = {tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533, tmp533};
    assign tmp535 = {tmp534, const_67_0};
    assign tmp536 = tmp13 - tmp535;
    assign tmp537 = {tmp536[256]};
    assign tmp538 = {tmp13[255]};
    assign tmp539 = ~tmp538;
    assign tmp540 = tmp537 ^ tmp539;
    assign tmp541 = {tmp535[255]};
    assign tmp542 = ~tmp541;
    assign tmp543 = tmp540 ^ tmp542;
    assign tmp544 = tmp531 & tmp543;
    assign tmp545 = {const_68_0};
    assign tmp546 = {tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545, tmp545};
    assign tmp547 = {tmp546, const_68_0};
    assign tmp548 = {tmp479[255]};
    assign tmp549 = tmp547 - tmp479;
    assign tmp550 = {tmp549[256]};
    assign tmp551 = {tmp547[255]};
    assign tmp552 = ~tmp551;
    assign tmp553 = tmp550 ^ tmp552;
    assign tmp554 = {tmp479[255]};
    assign tmp555 = ~tmp554;
    assign tmp556 = tmp553 ^ tmp555;
    assign tmp557 = tmp547 == tmp479;
    assign tmp558 = tmp556 | tmp557;
    assign tmp559 = tmp544 & tmp558;
    assign tmp560 = tmp519 ? const_69_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp479;
    assign tmp561 = tmp559 ? _ver_out_tmp_30 : tmp560;
    assign tmp562 = ~tmp35;
    assign tmp563 = ~tmp36;
    assign tmp564 = tmp562 & tmp563;
    assign tmp565 = tmp564 & tmp57;
    assign tmp566 = ~tmp68;
    assign tmp567 = tmp565 & tmp566;
    assign tmp568 = ~tmp69;
    assign tmp569 = tmp567 & tmp568;
    assign tmp570 = ~tmp108;
    assign tmp571 = tmp569 & tmp570;
    assign tmp572 = ~tmp375;
    assign tmp573 = tmp571 & tmp572;
    assign tmp574 = tmp573 & tmp470;
    assign tmp575 = ~tmp35;
    assign tmp576 = ~tmp36;
    assign tmp577 = tmp575 & tmp576;
    assign tmp578 = tmp577 & tmp57;
    assign tmp579 = ~tmp68;
    assign tmp580 = tmp578 & tmp579;
    assign tmp581 = ~tmp69;
    assign tmp582 = tmp580 & tmp581;
    assign tmp583 = ~tmp108;
    assign tmp584 = tmp582 & tmp583;
    assign tmp585 = ~tmp375;
    assign tmp586 = tmp584 & tmp585;
    assign tmp587 = tmp586 & tmp470;
    assign tmp588 = {tmp12[255]};
    assign tmp589 = {tmp588};
    assign tmp590 = {tmp589, tmp12};
    assign tmp591 = {tmp14[255]};
    assign tmp592 = {tmp591};
    assign tmp593 = {tmp592, tmp14};
    assign tmp594 = tmp590 + tmp593;
    assign tmp595 = {tmp594[256], tmp594[255], tmp594[254], tmp594[253], tmp594[252], tmp594[251], tmp594[250], tmp594[249], tmp594[248], tmp594[247], tmp594[246], tmp594[245], tmp594[244], tmp594[243], tmp594[242], tmp594[241], tmp594[240], tmp594[239], tmp594[238], tmp594[237], tmp594[236], tmp594[235], tmp594[234], tmp594[233], tmp594[232], tmp594[231], tmp594[230], tmp594[229], tmp594[228], tmp594[227], tmp594[226], tmp594[225], tmp594[224], tmp594[223], tmp594[222], tmp594[221], tmp594[220], tmp594[219], tmp594[218], tmp594[217], tmp594[216], tmp594[215], tmp594[214], tmp594[213], tmp594[212], tmp594[211], tmp594[210], tmp594[209], tmp594[208], tmp594[207], tmp594[206], tmp594[205], tmp594[204], tmp594[203], tmp594[202], tmp594[201], tmp594[200], tmp594[199], tmp594[198], tmp594[197], tmp594[196], tmp594[195], tmp594[194], tmp594[193], tmp594[192], tmp594[191], tmp594[190], tmp594[189], tmp594[188], tmp594[187], tmp594[186], tmp594[185], tmp594[184], tmp594[183], tmp594[182], tmp594[181], tmp594[180], tmp594[179], tmp594[178], tmp594[177], tmp594[176], tmp594[175], tmp594[174], tmp594[173], tmp594[172], tmp594[171], tmp594[170], tmp594[169], tmp594[168], tmp594[167], tmp594[166], tmp594[165], tmp594[164], tmp594[163], tmp594[162], tmp594[161], tmp594[160], tmp594[159], tmp594[158], tmp594[157], tmp594[156], tmp594[155], tmp594[154], tmp594[153], tmp594[152], tmp594[151], tmp594[150], tmp594[149], tmp594[148], tmp594[147], tmp594[146], tmp594[145], tmp594[144], tmp594[143], tmp594[142], tmp594[141], tmp594[140], tmp594[139], tmp594[138], tmp594[137], tmp594[136], tmp594[135], tmp594[134], tmp594[133], tmp594[132], tmp594[131], tmp594[130], tmp594[129], tmp594[128], tmp594[127], tmp594[126], tmp594[125], tmp594[124], tmp594[123], tmp594[122], tmp594[121], tmp594[120], tmp594[119], tmp594[118], tmp594[117], tmp594[116], tmp594[115], tmp594[114], tmp594[113], tmp594[112], tmp594[111], tmp594[110], tmp594[109], tmp594[108], tmp594[107], tmp594[106], tmp594[105], tmp594[104], tmp594[103], tmp594[102], tmp594[101], tmp594[100], tmp594[99], tmp594[98], tmp594[97], tmp594[96], tmp594[95], tmp594[94], tmp594[93], tmp594[92], tmp594[91], tmp594[90], tmp594[89], tmp594[88], tmp594[87], tmp594[86], tmp594[85], tmp594[84], tmp594[83], tmp594[82], tmp594[81], tmp594[80], tmp594[79], tmp594[78], tmp594[77], tmp594[76], tmp594[75], tmp594[74], tmp594[73], tmp594[72], tmp594[71], tmp594[70], tmp594[69], tmp594[68], tmp594[67], tmp594[66], tmp594[65], tmp594[64], tmp594[63], tmp594[62], tmp594[61], tmp594[60], tmp594[59], tmp594[58], tmp594[57], tmp594[56], tmp594[55], tmp594[54], tmp594[53], tmp594[52], tmp594[51], tmp594[50], tmp594[49], tmp594[48], tmp594[47], tmp594[46], tmp594[45], tmp594[44], tmp594[43], tmp594[42], tmp594[41], tmp594[40], tmp594[39], tmp594[38], tmp594[37], tmp594[36], tmp594[35], tmp594[34], tmp594[33], tmp594[32], tmp594[31], tmp594[30], tmp594[29], tmp594[28], tmp594[27], tmp594[26], tmp594[25], tmp594[24], tmp594[23], tmp594[22], tmp594[21], tmp594[20], tmp594[19], tmp594[18], tmp594[17], tmp594[16], tmp594[15], tmp594[14], tmp594[13], tmp594[12], tmp594[11], tmp594[10], tmp594[9], tmp594[8], tmp594[7], tmp594[6], tmp594[5], tmp594[4], tmp594[3], tmp594[2], tmp594[1], tmp594[0]};
    assign tmp596 = {tmp595[255], tmp595[254], tmp595[253], tmp595[252], tmp595[251], tmp595[250], tmp595[249], tmp595[248], tmp595[247], tmp595[246], tmp595[245], tmp595[244], tmp595[243], tmp595[242], tmp595[241], tmp595[240], tmp595[239], tmp595[238], tmp595[237], tmp595[236], tmp595[235], tmp595[234], tmp595[233], tmp595[232], tmp595[231], tmp595[230], tmp595[229], tmp595[228], tmp595[227], tmp595[226], tmp595[225], tmp595[224], tmp595[223], tmp595[222], tmp595[221], tmp595[220], tmp595[219], tmp595[218], tmp595[217], tmp595[216], tmp595[215], tmp595[214], tmp595[213], tmp595[212], tmp595[211], tmp595[210], tmp595[209], tmp595[208], tmp595[207], tmp595[206], tmp595[205], tmp595[204], tmp595[203], tmp595[202], tmp595[201], tmp595[200], tmp595[199], tmp595[198], tmp595[197], tmp595[196], tmp595[195], tmp595[194], tmp595[193], tmp595[192], tmp595[191], tmp595[190], tmp595[189], tmp595[188], tmp595[187], tmp595[186], tmp595[185], tmp595[184], tmp595[183], tmp595[182], tmp595[181], tmp595[180], tmp595[179], tmp595[178], tmp595[177], tmp595[176], tmp595[175], tmp595[174], tmp595[173], tmp595[172], tmp595[171], tmp595[170], tmp595[169], tmp595[168], tmp595[167], tmp595[166], tmp595[165], tmp595[164], tmp595[163], tmp595[162], tmp595[161], tmp595[160], tmp595[159], tmp595[158], tmp595[157], tmp595[156], tmp595[155], tmp595[154], tmp595[153], tmp595[152], tmp595[151], tmp595[150], tmp595[149], tmp595[148], tmp595[147], tmp595[146], tmp595[145], tmp595[144], tmp595[143], tmp595[142], tmp595[141], tmp595[140], tmp595[139], tmp595[138], tmp595[137], tmp595[136], tmp595[135], tmp595[134], tmp595[133], tmp595[132], tmp595[131], tmp595[130], tmp595[129], tmp595[128], tmp595[127], tmp595[126], tmp595[125], tmp595[124], tmp595[123], tmp595[122], tmp595[121], tmp595[120], tmp595[119], tmp595[118], tmp595[117], tmp595[116], tmp595[115], tmp595[114], tmp595[113], tmp595[112], tmp595[111], tmp595[110], tmp595[109], tmp595[108], tmp595[107], tmp595[106], tmp595[105], tmp595[104], tmp595[103], tmp595[102], tmp595[101], tmp595[100], tmp595[99], tmp595[98], tmp595[97], tmp595[96], tmp595[95], tmp595[94], tmp595[93], tmp595[92], tmp595[91], tmp595[90], tmp595[89], tmp595[88], tmp595[87], tmp595[86], tmp595[85], tmp595[84], tmp595[83], tmp595[82], tmp595[81], tmp595[80], tmp595[79], tmp595[78], tmp595[77], tmp595[76], tmp595[75], tmp595[74], tmp595[73], tmp595[72], tmp595[71], tmp595[70], tmp595[69], tmp595[68], tmp595[67], tmp595[66], tmp595[65], tmp595[64], tmp595[63], tmp595[62], tmp595[61], tmp595[60], tmp595[59], tmp595[58], tmp595[57], tmp595[56], tmp595[55], tmp595[54], tmp595[53], tmp595[52], tmp595[51], tmp595[50], tmp595[49], tmp595[48], tmp595[47], tmp595[46], tmp595[45], tmp595[44], tmp595[43], tmp595[42], tmp595[41], tmp595[40], tmp595[39], tmp595[38], tmp595[37], tmp595[36], tmp595[35], tmp595[34], tmp595[33], tmp595[32], tmp595[31], tmp595[30], tmp595[29], tmp595[28], tmp595[27], tmp595[26], tmp595[25], tmp595[24], tmp595[23], tmp595[22], tmp595[21], tmp595[20], tmp595[19], tmp595[18], tmp595[17], tmp595[16], tmp595[15], tmp595[14], tmp595[13], tmp595[12], tmp595[11], tmp595[10], tmp595[9], tmp595[8], tmp595[7], tmp595[6], tmp595[5], tmp595[4], tmp595[3], tmp595[2], tmp595[1], tmp595[0]};
    assign tmp597 = {const_71_0};
    assign tmp598 = {tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597, tmp597};
    assign tmp599 = {tmp598, const_71_0};
    assign tmp600 = {tmp12[255]};
    assign tmp601 = tmp599 - tmp12;
    assign tmp602 = {tmp601[256]};
    assign tmp603 = {tmp599[255]};
    assign tmp604 = ~tmp603;
    assign tmp605 = tmp602 ^ tmp604;
    assign tmp606 = {tmp12[255]};
    assign tmp607 = ~tmp606;
    assign tmp608 = tmp605 ^ tmp607;
    assign tmp609 = {const_72_0};
    assign tmp610 = {tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609, tmp609};
    assign tmp611 = {tmp610, const_72_0};
    assign tmp612 = {tmp14[255]};
    assign tmp613 = tmp611 - tmp14;
    assign tmp614 = {tmp613[256]};
    assign tmp615 = {tmp611[255]};
    assign tmp616 = ~tmp615;
    assign tmp617 = tmp614 ^ tmp616;
    assign tmp618 = {tmp14[255]};
    assign tmp619 = ~tmp618;
    assign tmp620 = tmp617 ^ tmp619;
    assign tmp621 = tmp608 & tmp620;
    assign tmp622 = {tmp596[255]};
    assign tmp623 = {const_73_0};
    assign tmp624 = {tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623, tmp623};
    assign tmp625 = {tmp624, const_73_0};
    assign tmp626 = tmp596 - tmp625;
    assign tmp627 = {tmp626[256]};
    assign tmp628 = {tmp596[255]};
    assign tmp629 = ~tmp628;
    assign tmp630 = tmp627 ^ tmp629;
    assign tmp631 = {tmp625[255]};
    assign tmp632 = ~tmp631;
    assign tmp633 = tmp630 ^ tmp632;
    assign tmp634 = tmp596 == tmp625;
    assign tmp635 = tmp633 | tmp634;
    assign tmp636 = tmp621 & tmp635;
    assign tmp637 = {tmp12[255]};
    assign tmp638 = {const_74_0};
    assign tmp639 = {tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638, tmp638};
    assign tmp640 = {tmp639, const_74_0};
    assign tmp641 = tmp12 - tmp640;
    assign tmp642 = {tmp641[256]};
    assign tmp643 = {tmp12[255]};
    assign tmp644 = ~tmp643;
    assign tmp645 = tmp642 ^ tmp644;
    assign tmp646 = {tmp640[255]};
    assign tmp647 = ~tmp646;
    assign tmp648 = tmp645 ^ tmp647;
    assign tmp649 = {tmp14[255]};
    assign tmp650 = {const_75_0};
    assign tmp651 = {tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650, tmp650};
    assign tmp652 = {tmp651, const_75_0};
    assign tmp653 = tmp14 - tmp652;
    assign tmp654 = {tmp653[256]};
    assign tmp655 = {tmp14[255]};
    assign tmp656 = ~tmp655;
    assign tmp657 = tmp654 ^ tmp656;
    assign tmp658 = {tmp652[255]};
    assign tmp659 = ~tmp658;
    assign tmp660 = tmp657 ^ tmp659;
    assign tmp661 = tmp648 & tmp660;
    assign tmp662 = {const_76_0};
    assign tmp663 = {tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662, tmp662};
    assign tmp664 = {tmp663, const_76_0};
    assign tmp665 = {tmp596[255]};
    assign tmp666 = tmp664 - tmp596;
    assign tmp667 = {tmp666[256]};
    assign tmp668 = {tmp664[255]};
    assign tmp669 = ~tmp668;
    assign tmp670 = tmp667 ^ tmp669;
    assign tmp671 = {tmp596[255]};
    assign tmp672 = ~tmp671;
    assign tmp673 = tmp670 ^ tmp672;
    assign tmp674 = tmp664 == tmp596;
    assign tmp675 = tmp673 | tmp674;
    assign tmp676 = tmp661 & tmp675;
    assign tmp677 = tmp636 ? const_77_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp596;
    assign tmp678 = tmp676 ? _ver_out_tmp_33 : tmp677;
    assign tmp679 = ~tmp35;
    assign tmp680 = ~tmp36;
    assign tmp681 = tmp679 & tmp680;
    assign tmp682 = tmp681 & tmp57;
    assign tmp683 = ~tmp68;
    assign tmp684 = tmp682 & tmp683;
    assign tmp685 = ~tmp69;
    assign tmp686 = tmp684 & tmp685;
    assign tmp687 = ~tmp108;
    assign tmp688 = tmp686 & tmp687;
    assign tmp689 = ~tmp375;
    assign tmp690 = tmp688 & tmp689;
    assign tmp691 = tmp690 & tmp470;
    assign tmp692 = ~tmp35;
    assign tmp693 = ~tmp36;
    assign tmp694 = tmp692 & tmp693;
    assign tmp695 = tmp694 & tmp57;
    assign tmp696 = ~tmp68;
    assign tmp697 = tmp695 & tmp696;
    assign tmp698 = ~tmp69;
    assign tmp699 = tmp697 & tmp698;
    assign tmp700 = ~tmp108;
    assign tmp701 = tmp699 & tmp700;
    assign tmp702 = ~tmp375;
    assign tmp703 = tmp701 & tmp702;
    assign tmp704 = tmp703 & tmp470;
    assign tmp705 = {tmp15[255]};
    assign tmp706 = {tmp705};
    assign tmp707 = {tmp706, tmp15};
    assign tmp708 = {tmp17[255]};
    assign tmp709 = {tmp708};
    assign tmp710 = {tmp709, tmp17};
    assign tmp711 = tmp707 + tmp710;
    assign tmp712 = {tmp711[256], tmp711[255], tmp711[254], tmp711[253], tmp711[252], tmp711[251], tmp711[250], tmp711[249], tmp711[248], tmp711[247], tmp711[246], tmp711[245], tmp711[244], tmp711[243], tmp711[242], tmp711[241], tmp711[240], tmp711[239], tmp711[238], tmp711[237], tmp711[236], tmp711[235], tmp711[234], tmp711[233], tmp711[232], tmp711[231], tmp711[230], tmp711[229], tmp711[228], tmp711[227], tmp711[226], tmp711[225], tmp711[224], tmp711[223], tmp711[222], tmp711[221], tmp711[220], tmp711[219], tmp711[218], tmp711[217], tmp711[216], tmp711[215], tmp711[214], tmp711[213], tmp711[212], tmp711[211], tmp711[210], tmp711[209], tmp711[208], tmp711[207], tmp711[206], tmp711[205], tmp711[204], tmp711[203], tmp711[202], tmp711[201], tmp711[200], tmp711[199], tmp711[198], tmp711[197], tmp711[196], tmp711[195], tmp711[194], tmp711[193], tmp711[192], tmp711[191], tmp711[190], tmp711[189], tmp711[188], tmp711[187], tmp711[186], tmp711[185], tmp711[184], tmp711[183], tmp711[182], tmp711[181], tmp711[180], tmp711[179], tmp711[178], tmp711[177], tmp711[176], tmp711[175], tmp711[174], tmp711[173], tmp711[172], tmp711[171], tmp711[170], tmp711[169], tmp711[168], tmp711[167], tmp711[166], tmp711[165], tmp711[164], tmp711[163], tmp711[162], tmp711[161], tmp711[160], tmp711[159], tmp711[158], tmp711[157], tmp711[156], tmp711[155], tmp711[154], tmp711[153], tmp711[152], tmp711[151], tmp711[150], tmp711[149], tmp711[148], tmp711[147], tmp711[146], tmp711[145], tmp711[144], tmp711[143], tmp711[142], tmp711[141], tmp711[140], tmp711[139], tmp711[138], tmp711[137], tmp711[136], tmp711[135], tmp711[134], tmp711[133], tmp711[132], tmp711[131], tmp711[130], tmp711[129], tmp711[128], tmp711[127], tmp711[126], tmp711[125], tmp711[124], tmp711[123], tmp711[122], tmp711[121], tmp711[120], tmp711[119], tmp711[118], tmp711[117], tmp711[116], tmp711[115], tmp711[114], tmp711[113], tmp711[112], tmp711[111], tmp711[110], tmp711[109], tmp711[108], tmp711[107], tmp711[106], tmp711[105], tmp711[104], tmp711[103], tmp711[102], tmp711[101], tmp711[100], tmp711[99], tmp711[98], tmp711[97], tmp711[96], tmp711[95], tmp711[94], tmp711[93], tmp711[92], tmp711[91], tmp711[90], tmp711[89], tmp711[88], tmp711[87], tmp711[86], tmp711[85], tmp711[84], tmp711[83], tmp711[82], tmp711[81], tmp711[80], tmp711[79], tmp711[78], tmp711[77], tmp711[76], tmp711[75], tmp711[74], tmp711[73], tmp711[72], tmp711[71], tmp711[70], tmp711[69], tmp711[68], tmp711[67], tmp711[66], tmp711[65], tmp711[64], tmp711[63], tmp711[62], tmp711[61], tmp711[60], tmp711[59], tmp711[58], tmp711[57], tmp711[56], tmp711[55], tmp711[54], tmp711[53], tmp711[52], tmp711[51], tmp711[50], tmp711[49], tmp711[48], tmp711[47], tmp711[46], tmp711[45], tmp711[44], tmp711[43], tmp711[42], tmp711[41], tmp711[40], tmp711[39], tmp711[38], tmp711[37], tmp711[36], tmp711[35], tmp711[34], tmp711[33], tmp711[32], tmp711[31], tmp711[30], tmp711[29], tmp711[28], tmp711[27], tmp711[26], tmp711[25], tmp711[24], tmp711[23], tmp711[22], tmp711[21], tmp711[20], tmp711[19], tmp711[18], tmp711[17], tmp711[16], tmp711[15], tmp711[14], tmp711[13], tmp711[12], tmp711[11], tmp711[10], tmp711[9], tmp711[8], tmp711[7], tmp711[6], tmp711[5], tmp711[4], tmp711[3], tmp711[2], tmp711[1], tmp711[0]};
    assign tmp713 = {tmp712[255], tmp712[254], tmp712[253], tmp712[252], tmp712[251], tmp712[250], tmp712[249], tmp712[248], tmp712[247], tmp712[246], tmp712[245], tmp712[244], tmp712[243], tmp712[242], tmp712[241], tmp712[240], tmp712[239], tmp712[238], tmp712[237], tmp712[236], tmp712[235], tmp712[234], tmp712[233], tmp712[232], tmp712[231], tmp712[230], tmp712[229], tmp712[228], tmp712[227], tmp712[226], tmp712[225], tmp712[224], tmp712[223], tmp712[222], tmp712[221], tmp712[220], tmp712[219], tmp712[218], tmp712[217], tmp712[216], tmp712[215], tmp712[214], tmp712[213], tmp712[212], tmp712[211], tmp712[210], tmp712[209], tmp712[208], tmp712[207], tmp712[206], tmp712[205], tmp712[204], tmp712[203], tmp712[202], tmp712[201], tmp712[200], tmp712[199], tmp712[198], tmp712[197], tmp712[196], tmp712[195], tmp712[194], tmp712[193], tmp712[192], tmp712[191], tmp712[190], tmp712[189], tmp712[188], tmp712[187], tmp712[186], tmp712[185], tmp712[184], tmp712[183], tmp712[182], tmp712[181], tmp712[180], tmp712[179], tmp712[178], tmp712[177], tmp712[176], tmp712[175], tmp712[174], tmp712[173], tmp712[172], tmp712[171], tmp712[170], tmp712[169], tmp712[168], tmp712[167], tmp712[166], tmp712[165], tmp712[164], tmp712[163], tmp712[162], tmp712[161], tmp712[160], tmp712[159], tmp712[158], tmp712[157], tmp712[156], tmp712[155], tmp712[154], tmp712[153], tmp712[152], tmp712[151], tmp712[150], tmp712[149], tmp712[148], tmp712[147], tmp712[146], tmp712[145], tmp712[144], tmp712[143], tmp712[142], tmp712[141], tmp712[140], tmp712[139], tmp712[138], tmp712[137], tmp712[136], tmp712[135], tmp712[134], tmp712[133], tmp712[132], tmp712[131], tmp712[130], tmp712[129], tmp712[128], tmp712[127], tmp712[126], tmp712[125], tmp712[124], tmp712[123], tmp712[122], tmp712[121], tmp712[120], tmp712[119], tmp712[118], tmp712[117], tmp712[116], tmp712[115], tmp712[114], tmp712[113], tmp712[112], tmp712[111], tmp712[110], tmp712[109], tmp712[108], tmp712[107], tmp712[106], tmp712[105], tmp712[104], tmp712[103], tmp712[102], tmp712[101], tmp712[100], tmp712[99], tmp712[98], tmp712[97], tmp712[96], tmp712[95], tmp712[94], tmp712[93], tmp712[92], tmp712[91], tmp712[90], tmp712[89], tmp712[88], tmp712[87], tmp712[86], tmp712[85], tmp712[84], tmp712[83], tmp712[82], tmp712[81], tmp712[80], tmp712[79], tmp712[78], tmp712[77], tmp712[76], tmp712[75], tmp712[74], tmp712[73], tmp712[72], tmp712[71], tmp712[70], tmp712[69], tmp712[68], tmp712[67], tmp712[66], tmp712[65], tmp712[64], tmp712[63], tmp712[62], tmp712[61], tmp712[60], tmp712[59], tmp712[58], tmp712[57], tmp712[56], tmp712[55], tmp712[54], tmp712[53], tmp712[52], tmp712[51], tmp712[50], tmp712[49], tmp712[48], tmp712[47], tmp712[46], tmp712[45], tmp712[44], tmp712[43], tmp712[42], tmp712[41], tmp712[40], tmp712[39], tmp712[38], tmp712[37], tmp712[36], tmp712[35], tmp712[34], tmp712[33], tmp712[32], tmp712[31], tmp712[30], tmp712[29], tmp712[28], tmp712[27], tmp712[26], tmp712[25], tmp712[24], tmp712[23], tmp712[22], tmp712[21], tmp712[20], tmp712[19], tmp712[18], tmp712[17], tmp712[16], tmp712[15], tmp712[14], tmp712[13], tmp712[12], tmp712[11], tmp712[10], tmp712[9], tmp712[8], tmp712[7], tmp712[6], tmp712[5], tmp712[4], tmp712[3], tmp712[2], tmp712[1], tmp712[0]};
    assign tmp714 = {const_79_0};
    assign tmp715 = {tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714, tmp714};
    assign tmp716 = {tmp715, const_79_0};
    assign tmp717 = {tmp15[255]};
    assign tmp718 = tmp716 - tmp15;
    assign tmp719 = {tmp718[256]};
    assign tmp720 = {tmp716[255]};
    assign tmp721 = ~tmp720;
    assign tmp722 = tmp719 ^ tmp721;
    assign tmp723 = {tmp15[255]};
    assign tmp724 = ~tmp723;
    assign tmp725 = tmp722 ^ tmp724;
    assign tmp726 = {const_80_0};
    assign tmp727 = {tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726, tmp726};
    assign tmp728 = {tmp727, const_80_0};
    assign tmp729 = {tmp17[255]};
    assign tmp730 = tmp728 - tmp17;
    assign tmp731 = {tmp730[256]};
    assign tmp732 = {tmp728[255]};
    assign tmp733 = ~tmp732;
    assign tmp734 = tmp731 ^ tmp733;
    assign tmp735 = {tmp17[255]};
    assign tmp736 = ~tmp735;
    assign tmp737 = tmp734 ^ tmp736;
    assign tmp738 = tmp725 & tmp737;
    assign tmp739 = {tmp713[255]};
    assign tmp740 = {const_81_0};
    assign tmp741 = {tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740, tmp740};
    assign tmp742 = {tmp741, const_81_0};
    assign tmp743 = tmp713 - tmp742;
    assign tmp744 = {tmp743[256]};
    assign tmp745 = {tmp713[255]};
    assign tmp746 = ~tmp745;
    assign tmp747 = tmp744 ^ tmp746;
    assign tmp748 = {tmp742[255]};
    assign tmp749 = ~tmp748;
    assign tmp750 = tmp747 ^ tmp749;
    assign tmp751 = tmp713 == tmp742;
    assign tmp752 = tmp750 | tmp751;
    assign tmp753 = tmp738 & tmp752;
    assign tmp754 = {tmp15[255]};
    assign tmp755 = {const_82_0};
    assign tmp756 = {tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755, tmp755};
    assign tmp757 = {tmp756, const_82_0};
    assign tmp758 = tmp15 - tmp757;
    assign tmp759 = {tmp758[256]};
    assign tmp760 = {tmp15[255]};
    assign tmp761 = ~tmp760;
    assign tmp762 = tmp759 ^ tmp761;
    assign tmp763 = {tmp757[255]};
    assign tmp764 = ~tmp763;
    assign tmp765 = tmp762 ^ tmp764;
    assign tmp766 = {tmp17[255]};
    assign tmp767 = {const_83_0};
    assign tmp768 = {tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767, tmp767};
    assign tmp769 = {tmp768, const_83_0};
    assign tmp770 = tmp17 - tmp769;
    assign tmp771 = {tmp770[256]};
    assign tmp772 = {tmp17[255]};
    assign tmp773 = ~tmp772;
    assign tmp774 = tmp771 ^ tmp773;
    assign tmp775 = {tmp769[255]};
    assign tmp776 = ~tmp775;
    assign tmp777 = tmp774 ^ tmp776;
    assign tmp778 = tmp765 & tmp777;
    assign tmp779 = {const_84_0};
    assign tmp780 = {tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779, tmp779};
    assign tmp781 = {tmp780, const_84_0};
    assign tmp782 = {tmp713[255]};
    assign tmp783 = tmp781 - tmp713;
    assign tmp784 = {tmp783[256]};
    assign tmp785 = {tmp781[255]};
    assign tmp786 = ~tmp785;
    assign tmp787 = tmp784 ^ tmp786;
    assign tmp788 = {tmp713[255]};
    assign tmp789 = ~tmp788;
    assign tmp790 = tmp787 ^ tmp789;
    assign tmp791 = tmp781 == tmp713;
    assign tmp792 = tmp790 | tmp791;
    assign tmp793 = tmp778 & tmp792;
    assign tmp794 = tmp753 ? const_85_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp713;
    assign tmp795 = tmp793 ? _ver_out_tmp_38 : tmp794;
    assign tmp796 = ~tmp35;
    assign tmp797 = ~tmp36;
    assign tmp798 = tmp796 & tmp797;
    assign tmp799 = tmp798 & tmp57;
    assign tmp800 = ~tmp68;
    assign tmp801 = tmp799 & tmp800;
    assign tmp802 = ~tmp69;
    assign tmp803 = tmp801 & tmp802;
    assign tmp804 = ~tmp108;
    assign tmp805 = tmp803 & tmp804;
    assign tmp806 = ~tmp375;
    assign tmp807 = tmp805 & tmp806;
    assign tmp808 = tmp807 & tmp470;
    assign tmp809 = ~tmp35;
    assign tmp810 = ~tmp36;
    assign tmp811 = tmp809 & tmp810;
    assign tmp812 = tmp811 & tmp57;
    assign tmp813 = ~tmp68;
    assign tmp814 = tmp812 & tmp813;
    assign tmp815 = ~tmp69;
    assign tmp816 = tmp814 & tmp815;
    assign tmp817 = ~tmp108;
    assign tmp818 = tmp816 & tmp817;
    assign tmp819 = ~tmp375;
    assign tmp820 = tmp818 & tmp819;
    assign tmp821 = tmp820 & tmp470;
    assign tmp822 = {tmp16[255]};
    assign tmp823 = {tmp822};
    assign tmp824 = {tmp823, tmp16};
    assign tmp825 = {tmp18[255]};
    assign tmp826 = {tmp825};
    assign tmp827 = {tmp826, tmp18};
    assign tmp828 = tmp824 + tmp827;
    assign tmp829 = {tmp828[256], tmp828[255], tmp828[254], tmp828[253], tmp828[252], tmp828[251], tmp828[250], tmp828[249], tmp828[248], tmp828[247], tmp828[246], tmp828[245], tmp828[244], tmp828[243], tmp828[242], tmp828[241], tmp828[240], tmp828[239], tmp828[238], tmp828[237], tmp828[236], tmp828[235], tmp828[234], tmp828[233], tmp828[232], tmp828[231], tmp828[230], tmp828[229], tmp828[228], tmp828[227], tmp828[226], tmp828[225], tmp828[224], tmp828[223], tmp828[222], tmp828[221], tmp828[220], tmp828[219], tmp828[218], tmp828[217], tmp828[216], tmp828[215], tmp828[214], tmp828[213], tmp828[212], tmp828[211], tmp828[210], tmp828[209], tmp828[208], tmp828[207], tmp828[206], tmp828[205], tmp828[204], tmp828[203], tmp828[202], tmp828[201], tmp828[200], tmp828[199], tmp828[198], tmp828[197], tmp828[196], tmp828[195], tmp828[194], tmp828[193], tmp828[192], tmp828[191], tmp828[190], tmp828[189], tmp828[188], tmp828[187], tmp828[186], tmp828[185], tmp828[184], tmp828[183], tmp828[182], tmp828[181], tmp828[180], tmp828[179], tmp828[178], tmp828[177], tmp828[176], tmp828[175], tmp828[174], tmp828[173], tmp828[172], tmp828[171], tmp828[170], tmp828[169], tmp828[168], tmp828[167], tmp828[166], tmp828[165], tmp828[164], tmp828[163], tmp828[162], tmp828[161], tmp828[160], tmp828[159], tmp828[158], tmp828[157], tmp828[156], tmp828[155], tmp828[154], tmp828[153], tmp828[152], tmp828[151], tmp828[150], tmp828[149], tmp828[148], tmp828[147], tmp828[146], tmp828[145], tmp828[144], tmp828[143], tmp828[142], tmp828[141], tmp828[140], tmp828[139], tmp828[138], tmp828[137], tmp828[136], tmp828[135], tmp828[134], tmp828[133], tmp828[132], tmp828[131], tmp828[130], tmp828[129], tmp828[128], tmp828[127], tmp828[126], tmp828[125], tmp828[124], tmp828[123], tmp828[122], tmp828[121], tmp828[120], tmp828[119], tmp828[118], tmp828[117], tmp828[116], tmp828[115], tmp828[114], tmp828[113], tmp828[112], tmp828[111], tmp828[110], tmp828[109], tmp828[108], tmp828[107], tmp828[106], tmp828[105], tmp828[104], tmp828[103], tmp828[102], tmp828[101], tmp828[100], tmp828[99], tmp828[98], tmp828[97], tmp828[96], tmp828[95], tmp828[94], tmp828[93], tmp828[92], tmp828[91], tmp828[90], tmp828[89], tmp828[88], tmp828[87], tmp828[86], tmp828[85], tmp828[84], tmp828[83], tmp828[82], tmp828[81], tmp828[80], tmp828[79], tmp828[78], tmp828[77], tmp828[76], tmp828[75], tmp828[74], tmp828[73], tmp828[72], tmp828[71], tmp828[70], tmp828[69], tmp828[68], tmp828[67], tmp828[66], tmp828[65], tmp828[64], tmp828[63], tmp828[62], tmp828[61], tmp828[60], tmp828[59], tmp828[58], tmp828[57], tmp828[56], tmp828[55], tmp828[54], tmp828[53], tmp828[52], tmp828[51], tmp828[50], tmp828[49], tmp828[48], tmp828[47], tmp828[46], tmp828[45], tmp828[44], tmp828[43], tmp828[42], tmp828[41], tmp828[40], tmp828[39], tmp828[38], tmp828[37], tmp828[36], tmp828[35], tmp828[34], tmp828[33], tmp828[32], tmp828[31], tmp828[30], tmp828[29], tmp828[28], tmp828[27], tmp828[26], tmp828[25], tmp828[24], tmp828[23], tmp828[22], tmp828[21], tmp828[20], tmp828[19], tmp828[18], tmp828[17], tmp828[16], tmp828[15], tmp828[14], tmp828[13], tmp828[12], tmp828[11], tmp828[10], tmp828[9], tmp828[8], tmp828[7], tmp828[6], tmp828[5], tmp828[4], tmp828[3], tmp828[2], tmp828[1], tmp828[0]};
    assign tmp830 = {tmp829[255], tmp829[254], tmp829[253], tmp829[252], tmp829[251], tmp829[250], tmp829[249], tmp829[248], tmp829[247], tmp829[246], tmp829[245], tmp829[244], tmp829[243], tmp829[242], tmp829[241], tmp829[240], tmp829[239], tmp829[238], tmp829[237], tmp829[236], tmp829[235], tmp829[234], tmp829[233], tmp829[232], tmp829[231], tmp829[230], tmp829[229], tmp829[228], tmp829[227], tmp829[226], tmp829[225], tmp829[224], tmp829[223], tmp829[222], tmp829[221], tmp829[220], tmp829[219], tmp829[218], tmp829[217], tmp829[216], tmp829[215], tmp829[214], tmp829[213], tmp829[212], tmp829[211], tmp829[210], tmp829[209], tmp829[208], tmp829[207], tmp829[206], tmp829[205], tmp829[204], tmp829[203], tmp829[202], tmp829[201], tmp829[200], tmp829[199], tmp829[198], tmp829[197], tmp829[196], tmp829[195], tmp829[194], tmp829[193], tmp829[192], tmp829[191], tmp829[190], tmp829[189], tmp829[188], tmp829[187], tmp829[186], tmp829[185], tmp829[184], tmp829[183], tmp829[182], tmp829[181], tmp829[180], tmp829[179], tmp829[178], tmp829[177], tmp829[176], tmp829[175], tmp829[174], tmp829[173], tmp829[172], tmp829[171], tmp829[170], tmp829[169], tmp829[168], tmp829[167], tmp829[166], tmp829[165], tmp829[164], tmp829[163], tmp829[162], tmp829[161], tmp829[160], tmp829[159], tmp829[158], tmp829[157], tmp829[156], tmp829[155], tmp829[154], tmp829[153], tmp829[152], tmp829[151], tmp829[150], tmp829[149], tmp829[148], tmp829[147], tmp829[146], tmp829[145], tmp829[144], tmp829[143], tmp829[142], tmp829[141], tmp829[140], tmp829[139], tmp829[138], tmp829[137], tmp829[136], tmp829[135], tmp829[134], tmp829[133], tmp829[132], tmp829[131], tmp829[130], tmp829[129], tmp829[128], tmp829[127], tmp829[126], tmp829[125], tmp829[124], tmp829[123], tmp829[122], tmp829[121], tmp829[120], tmp829[119], tmp829[118], tmp829[117], tmp829[116], tmp829[115], tmp829[114], tmp829[113], tmp829[112], tmp829[111], tmp829[110], tmp829[109], tmp829[108], tmp829[107], tmp829[106], tmp829[105], tmp829[104], tmp829[103], tmp829[102], tmp829[101], tmp829[100], tmp829[99], tmp829[98], tmp829[97], tmp829[96], tmp829[95], tmp829[94], tmp829[93], tmp829[92], tmp829[91], tmp829[90], tmp829[89], tmp829[88], tmp829[87], tmp829[86], tmp829[85], tmp829[84], tmp829[83], tmp829[82], tmp829[81], tmp829[80], tmp829[79], tmp829[78], tmp829[77], tmp829[76], tmp829[75], tmp829[74], tmp829[73], tmp829[72], tmp829[71], tmp829[70], tmp829[69], tmp829[68], tmp829[67], tmp829[66], tmp829[65], tmp829[64], tmp829[63], tmp829[62], tmp829[61], tmp829[60], tmp829[59], tmp829[58], tmp829[57], tmp829[56], tmp829[55], tmp829[54], tmp829[53], tmp829[52], tmp829[51], tmp829[50], tmp829[49], tmp829[48], tmp829[47], tmp829[46], tmp829[45], tmp829[44], tmp829[43], tmp829[42], tmp829[41], tmp829[40], tmp829[39], tmp829[38], tmp829[37], tmp829[36], tmp829[35], tmp829[34], tmp829[33], tmp829[32], tmp829[31], tmp829[30], tmp829[29], tmp829[28], tmp829[27], tmp829[26], tmp829[25], tmp829[24], tmp829[23], tmp829[22], tmp829[21], tmp829[20], tmp829[19], tmp829[18], tmp829[17], tmp829[16], tmp829[15], tmp829[14], tmp829[13], tmp829[12], tmp829[11], tmp829[10], tmp829[9], tmp829[8], tmp829[7], tmp829[6], tmp829[5], tmp829[4], tmp829[3], tmp829[2], tmp829[1], tmp829[0]};
    assign tmp831 = {const_87_0};
    assign tmp832 = {tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831, tmp831};
    assign tmp833 = {tmp832, const_87_0};
    assign tmp834 = {tmp16[255]};
    assign tmp835 = tmp833 - tmp16;
    assign tmp836 = {tmp835[256]};
    assign tmp837 = {tmp833[255]};
    assign tmp838 = ~tmp837;
    assign tmp839 = tmp836 ^ tmp838;
    assign tmp840 = {tmp16[255]};
    assign tmp841 = ~tmp840;
    assign tmp842 = tmp839 ^ tmp841;
    assign tmp843 = {const_88_0};
    assign tmp844 = {tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843, tmp843};
    assign tmp845 = {tmp844, const_88_0};
    assign tmp846 = {tmp18[255]};
    assign tmp847 = tmp845 - tmp18;
    assign tmp848 = {tmp847[256]};
    assign tmp849 = {tmp845[255]};
    assign tmp850 = ~tmp849;
    assign tmp851 = tmp848 ^ tmp850;
    assign tmp852 = {tmp18[255]};
    assign tmp853 = ~tmp852;
    assign tmp854 = tmp851 ^ tmp853;
    assign tmp855 = tmp842 & tmp854;
    assign tmp856 = {tmp830[255]};
    assign tmp857 = {const_89_0};
    assign tmp858 = {tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857, tmp857};
    assign tmp859 = {tmp858, const_89_0};
    assign tmp860 = tmp830 - tmp859;
    assign tmp861 = {tmp860[256]};
    assign tmp862 = {tmp830[255]};
    assign tmp863 = ~tmp862;
    assign tmp864 = tmp861 ^ tmp863;
    assign tmp865 = {tmp859[255]};
    assign tmp866 = ~tmp865;
    assign tmp867 = tmp864 ^ tmp866;
    assign tmp868 = tmp830 == tmp859;
    assign tmp869 = tmp867 | tmp868;
    assign tmp870 = tmp855 & tmp869;
    assign tmp871 = {tmp16[255]};
    assign tmp872 = {const_90_0};
    assign tmp873 = {tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872, tmp872};
    assign tmp874 = {tmp873, const_90_0};
    assign tmp875 = tmp16 - tmp874;
    assign tmp876 = {tmp875[256]};
    assign tmp877 = {tmp16[255]};
    assign tmp878 = ~tmp877;
    assign tmp879 = tmp876 ^ tmp878;
    assign tmp880 = {tmp874[255]};
    assign tmp881 = ~tmp880;
    assign tmp882 = tmp879 ^ tmp881;
    assign tmp883 = {tmp18[255]};
    assign tmp884 = {const_91_0};
    assign tmp885 = {tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884, tmp884};
    assign tmp886 = {tmp885, const_91_0};
    assign tmp887 = tmp18 - tmp886;
    assign tmp888 = {tmp887[256]};
    assign tmp889 = {tmp18[255]};
    assign tmp890 = ~tmp889;
    assign tmp891 = tmp888 ^ tmp890;
    assign tmp892 = {tmp886[255]};
    assign tmp893 = ~tmp892;
    assign tmp894 = tmp891 ^ tmp893;
    assign tmp895 = tmp882 & tmp894;
    assign tmp896 = {const_92_0};
    assign tmp897 = {tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896, tmp896};
    assign tmp898 = {tmp897, const_92_0};
    assign tmp899 = {tmp830[255]};
    assign tmp900 = tmp898 - tmp830;
    assign tmp901 = {tmp900[256]};
    assign tmp902 = {tmp898[255]};
    assign tmp903 = ~tmp902;
    assign tmp904 = tmp901 ^ tmp903;
    assign tmp905 = {tmp830[255]};
    assign tmp906 = ~tmp905;
    assign tmp907 = tmp904 ^ tmp906;
    assign tmp908 = tmp898 == tmp830;
    assign tmp909 = tmp907 | tmp908;
    assign tmp910 = tmp895 & tmp909;
    assign tmp911 = tmp870 ? const_93_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp830;
    assign tmp912 = tmp910 ? _ver_out_tmp_40 : tmp911;
    assign tmp913 = ~tmp35;
    assign tmp914 = ~tmp36;
    assign tmp915 = tmp913 & tmp914;
    assign tmp916 = tmp915 & tmp57;
    assign tmp917 = ~tmp68;
    assign tmp918 = tmp916 & tmp917;
    assign tmp919 = ~tmp69;
    assign tmp920 = tmp918 & tmp919;
    assign tmp921 = ~tmp108;
    assign tmp922 = tmp920 & tmp921;
    assign tmp923 = ~tmp375;
    assign tmp924 = tmp922 & tmp923;
    assign tmp925 = tmp924 & tmp470;
    assign tmp926 = ~tmp35;
    assign tmp927 = ~tmp36;
    assign tmp928 = tmp926 & tmp927;
    assign tmp929 = tmp928 & tmp57;
    assign tmp930 = ~tmp68;
    assign tmp931 = tmp929 & tmp930;
    assign tmp932 = ~tmp69;
    assign tmp933 = tmp931 & tmp932;
    assign tmp934 = ~tmp108;
    assign tmp935 = tmp933 & tmp934;
    assign tmp936 = ~tmp375;
    assign tmp937 = tmp935 & tmp936;
    assign tmp938 = tmp937 & tmp470;
    assign tmp939 = my_calculator_in_x == const_95_8;
    assign tmp940 = tmp11 == _ver_out_tmp_41;
    assign tmp941 = {const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0, const_98_0};
    assign tmp942 = {tmp941, const_97_0};
    assign tmp943 = tmp942 - tmp11;
    assign tmp944 = {const_100_0, const_100_0};
    assign tmp945 = {tmp944, const_99_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp946 = tmp940 ? tmp945 : tmp943;
    assign tmp947 = {tmp946[255], tmp946[254], tmp946[253], tmp946[252], tmp946[251], tmp946[250], tmp946[249], tmp946[248], tmp946[247], tmp946[246], tmp946[245], tmp946[244], tmp946[243], tmp946[242], tmp946[241], tmp946[240], tmp946[239], tmp946[238], tmp946[237], tmp946[236], tmp946[235], tmp946[234], tmp946[233], tmp946[232], tmp946[231], tmp946[230], tmp946[229], tmp946[228], tmp946[227], tmp946[226], tmp946[225], tmp946[224], tmp946[223], tmp946[222], tmp946[221], tmp946[220], tmp946[219], tmp946[218], tmp946[217], tmp946[216], tmp946[215], tmp946[214], tmp946[213], tmp946[212], tmp946[211], tmp946[210], tmp946[209], tmp946[208], tmp946[207], tmp946[206], tmp946[205], tmp946[204], tmp946[203], tmp946[202], tmp946[201], tmp946[200], tmp946[199], tmp946[198], tmp946[197], tmp946[196], tmp946[195], tmp946[194], tmp946[193], tmp946[192], tmp946[191], tmp946[190], tmp946[189], tmp946[188], tmp946[187], tmp946[186], tmp946[185], tmp946[184], tmp946[183], tmp946[182], tmp946[181], tmp946[180], tmp946[179], tmp946[178], tmp946[177], tmp946[176], tmp946[175], tmp946[174], tmp946[173], tmp946[172], tmp946[171], tmp946[170], tmp946[169], tmp946[168], tmp946[167], tmp946[166], tmp946[165], tmp946[164], tmp946[163], tmp946[162], tmp946[161], tmp946[160], tmp946[159], tmp946[158], tmp946[157], tmp946[156], tmp946[155], tmp946[154], tmp946[153], tmp946[152], tmp946[151], tmp946[150], tmp946[149], tmp946[148], tmp946[147], tmp946[146], tmp946[145], tmp946[144], tmp946[143], tmp946[142], tmp946[141], tmp946[140], tmp946[139], tmp946[138], tmp946[137], tmp946[136], tmp946[135], tmp946[134], tmp946[133], tmp946[132], tmp946[131], tmp946[130], tmp946[129], tmp946[128], tmp946[127], tmp946[126], tmp946[125], tmp946[124], tmp946[123], tmp946[122], tmp946[121], tmp946[120], tmp946[119], tmp946[118], tmp946[117], tmp946[116], tmp946[115], tmp946[114], tmp946[113], tmp946[112], tmp946[111], tmp946[110], tmp946[109], tmp946[108], tmp946[107], tmp946[106], tmp946[105], tmp946[104], tmp946[103], tmp946[102], tmp946[101], tmp946[100], tmp946[99], tmp946[98], tmp946[97], tmp946[96], tmp946[95], tmp946[94], tmp946[93], tmp946[92], tmp946[91], tmp946[90], tmp946[89], tmp946[88], tmp946[87], tmp946[86], tmp946[85], tmp946[84], tmp946[83], tmp946[82], tmp946[81], tmp946[80], tmp946[79], tmp946[78], tmp946[77], tmp946[76], tmp946[75], tmp946[74], tmp946[73], tmp946[72], tmp946[71], tmp946[70], tmp946[69], tmp946[68], tmp946[67], tmp946[66], tmp946[65], tmp946[64], tmp946[63], tmp946[62], tmp946[61], tmp946[60], tmp946[59], tmp946[58], tmp946[57], tmp946[56], tmp946[55], tmp946[54], tmp946[53], tmp946[52], tmp946[51], tmp946[50], tmp946[49], tmp946[48], tmp946[47], tmp946[46], tmp946[45], tmp946[44], tmp946[43], tmp946[42], tmp946[41], tmp946[40], tmp946[39], tmp946[38], tmp946[37], tmp946[36], tmp946[35], tmp946[34], tmp946[33], tmp946[32], tmp946[31], tmp946[30], tmp946[29], tmp946[28], tmp946[27], tmp946[26], tmp946[25], tmp946[24], tmp946[23], tmp946[22], tmp946[21], tmp946[20], tmp946[19], tmp946[18], tmp946[17], tmp946[16], tmp946[15], tmp946[14], tmp946[13], tmp946[12], tmp946[11], tmp946[10], tmp946[9], tmp946[8], tmp946[7], tmp946[6], tmp946[5], tmp946[4], tmp946[3], tmp946[2], tmp946[1], tmp946[0]};
    assign tmp948 = ~tmp35;
    assign tmp949 = ~tmp36;
    assign tmp950 = tmp948 & tmp949;
    assign tmp951 = tmp950 & tmp57;
    assign tmp952 = ~tmp68;
    assign tmp953 = tmp951 & tmp952;
    assign tmp954 = ~tmp69;
    assign tmp955 = tmp953 & tmp954;
    assign tmp956 = ~tmp108;
    assign tmp957 = tmp955 & tmp956;
    assign tmp958 = ~tmp375;
    assign tmp959 = tmp957 & tmp958;
    assign tmp960 = ~tmp470;
    assign tmp961 = tmp959 & tmp960;
    assign tmp962 = tmp961 & tmp939;
    assign tmp963 = tmp12 == _ver_out_tmp_46;
    assign tmp964 = {const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0, const_103_0};
    assign tmp965 = {tmp964, const_102_0};
    assign tmp966 = tmp965 - tmp12;
    assign tmp967 = {const_105_0, const_105_0};
    assign tmp968 = {tmp967, const_104_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp969 = tmp963 ? tmp968 : tmp966;
    assign tmp970 = {tmp969[255], tmp969[254], tmp969[253], tmp969[252], tmp969[251], tmp969[250], tmp969[249], tmp969[248], tmp969[247], tmp969[246], tmp969[245], tmp969[244], tmp969[243], tmp969[242], tmp969[241], tmp969[240], tmp969[239], tmp969[238], tmp969[237], tmp969[236], tmp969[235], tmp969[234], tmp969[233], tmp969[232], tmp969[231], tmp969[230], tmp969[229], tmp969[228], tmp969[227], tmp969[226], tmp969[225], tmp969[224], tmp969[223], tmp969[222], tmp969[221], tmp969[220], tmp969[219], tmp969[218], tmp969[217], tmp969[216], tmp969[215], tmp969[214], tmp969[213], tmp969[212], tmp969[211], tmp969[210], tmp969[209], tmp969[208], tmp969[207], tmp969[206], tmp969[205], tmp969[204], tmp969[203], tmp969[202], tmp969[201], tmp969[200], tmp969[199], tmp969[198], tmp969[197], tmp969[196], tmp969[195], tmp969[194], tmp969[193], tmp969[192], tmp969[191], tmp969[190], tmp969[189], tmp969[188], tmp969[187], tmp969[186], tmp969[185], tmp969[184], tmp969[183], tmp969[182], tmp969[181], tmp969[180], tmp969[179], tmp969[178], tmp969[177], tmp969[176], tmp969[175], tmp969[174], tmp969[173], tmp969[172], tmp969[171], tmp969[170], tmp969[169], tmp969[168], tmp969[167], tmp969[166], tmp969[165], tmp969[164], tmp969[163], tmp969[162], tmp969[161], tmp969[160], tmp969[159], tmp969[158], tmp969[157], tmp969[156], tmp969[155], tmp969[154], tmp969[153], tmp969[152], tmp969[151], tmp969[150], tmp969[149], tmp969[148], tmp969[147], tmp969[146], tmp969[145], tmp969[144], tmp969[143], tmp969[142], tmp969[141], tmp969[140], tmp969[139], tmp969[138], tmp969[137], tmp969[136], tmp969[135], tmp969[134], tmp969[133], tmp969[132], tmp969[131], tmp969[130], tmp969[129], tmp969[128], tmp969[127], tmp969[126], tmp969[125], tmp969[124], tmp969[123], tmp969[122], tmp969[121], tmp969[120], tmp969[119], tmp969[118], tmp969[117], tmp969[116], tmp969[115], tmp969[114], tmp969[113], tmp969[112], tmp969[111], tmp969[110], tmp969[109], tmp969[108], tmp969[107], tmp969[106], tmp969[105], tmp969[104], tmp969[103], tmp969[102], tmp969[101], tmp969[100], tmp969[99], tmp969[98], tmp969[97], tmp969[96], tmp969[95], tmp969[94], tmp969[93], tmp969[92], tmp969[91], tmp969[90], tmp969[89], tmp969[88], tmp969[87], tmp969[86], tmp969[85], tmp969[84], tmp969[83], tmp969[82], tmp969[81], tmp969[80], tmp969[79], tmp969[78], tmp969[77], tmp969[76], tmp969[75], tmp969[74], tmp969[73], tmp969[72], tmp969[71], tmp969[70], tmp969[69], tmp969[68], tmp969[67], tmp969[66], tmp969[65], tmp969[64], tmp969[63], tmp969[62], tmp969[61], tmp969[60], tmp969[59], tmp969[58], tmp969[57], tmp969[56], tmp969[55], tmp969[54], tmp969[53], tmp969[52], tmp969[51], tmp969[50], tmp969[49], tmp969[48], tmp969[47], tmp969[46], tmp969[45], tmp969[44], tmp969[43], tmp969[42], tmp969[41], tmp969[40], tmp969[39], tmp969[38], tmp969[37], tmp969[36], tmp969[35], tmp969[34], tmp969[33], tmp969[32], tmp969[31], tmp969[30], tmp969[29], tmp969[28], tmp969[27], tmp969[26], tmp969[25], tmp969[24], tmp969[23], tmp969[22], tmp969[21], tmp969[20], tmp969[19], tmp969[18], tmp969[17], tmp969[16], tmp969[15], tmp969[14], tmp969[13], tmp969[12], tmp969[11], tmp969[10], tmp969[9], tmp969[8], tmp969[7], tmp969[6], tmp969[5], tmp969[4], tmp969[3], tmp969[2], tmp969[1], tmp969[0]};
    assign tmp971 = ~tmp35;
    assign tmp972 = ~tmp36;
    assign tmp973 = tmp971 & tmp972;
    assign tmp974 = tmp973 & tmp57;
    assign tmp975 = ~tmp68;
    assign tmp976 = tmp974 & tmp975;
    assign tmp977 = ~tmp69;
    assign tmp978 = tmp976 & tmp977;
    assign tmp979 = ~tmp108;
    assign tmp980 = tmp978 & tmp979;
    assign tmp981 = ~tmp375;
    assign tmp982 = tmp980 & tmp981;
    assign tmp983 = ~tmp470;
    assign tmp984 = tmp982 & tmp983;
    assign tmp985 = tmp984 & tmp939;
    assign tmp986 = tmp15 == _ver_out_tmp_48;
    assign tmp987 = {const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0, const_108_0};
    assign tmp988 = {tmp987, const_107_0};
    assign tmp989 = tmp988 - tmp15;
    assign tmp990 = {const_110_0, const_110_0};
    assign tmp991 = {tmp990, const_109_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp992 = tmp986 ? tmp991 : tmp989;
    assign tmp993 = {tmp992[255], tmp992[254], tmp992[253], tmp992[252], tmp992[251], tmp992[250], tmp992[249], tmp992[248], tmp992[247], tmp992[246], tmp992[245], tmp992[244], tmp992[243], tmp992[242], tmp992[241], tmp992[240], tmp992[239], tmp992[238], tmp992[237], tmp992[236], tmp992[235], tmp992[234], tmp992[233], tmp992[232], tmp992[231], tmp992[230], tmp992[229], tmp992[228], tmp992[227], tmp992[226], tmp992[225], tmp992[224], tmp992[223], tmp992[222], tmp992[221], tmp992[220], tmp992[219], tmp992[218], tmp992[217], tmp992[216], tmp992[215], tmp992[214], tmp992[213], tmp992[212], tmp992[211], tmp992[210], tmp992[209], tmp992[208], tmp992[207], tmp992[206], tmp992[205], tmp992[204], tmp992[203], tmp992[202], tmp992[201], tmp992[200], tmp992[199], tmp992[198], tmp992[197], tmp992[196], tmp992[195], tmp992[194], tmp992[193], tmp992[192], tmp992[191], tmp992[190], tmp992[189], tmp992[188], tmp992[187], tmp992[186], tmp992[185], tmp992[184], tmp992[183], tmp992[182], tmp992[181], tmp992[180], tmp992[179], tmp992[178], tmp992[177], tmp992[176], tmp992[175], tmp992[174], tmp992[173], tmp992[172], tmp992[171], tmp992[170], tmp992[169], tmp992[168], tmp992[167], tmp992[166], tmp992[165], tmp992[164], tmp992[163], tmp992[162], tmp992[161], tmp992[160], tmp992[159], tmp992[158], tmp992[157], tmp992[156], tmp992[155], tmp992[154], tmp992[153], tmp992[152], tmp992[151], tmp992[150], tmp992[149], tmp992[148], tmp992[147], tmp992[146], tmp992[145], tmp992[144], tmp992[143], tmp992[142], tmp992[141], tmp992[140], tmp992[139], tmp992[138], tmp992[137], tmp992[136], tmp992[135], tmp992[134], tmp992[133], tmp992[132], tmp992[131], tmp992[130], tmp992[129], tmp992[128], tmp992[127], tmp992[126], tmp992[125], tmp992[124], tmp992[123], tmp992[122], tmp992[121], tmp992[120], tmp992[119], tmp992[118], tmp992[117], tmp992[116], tmp992[115], tmp992[114], tmp992[113], tmp992[112], tmp992[111], tmp992[110], tmp992[109], tmp992[108], tmp992[107], tmp992[106], tmp992[105], tmp992[104], tmp992[103], tmp992[102], tmp992[101], tmp992[100], tmp992[99], tmp992[98], tmp992[97], tmp992[96], tmp992[95], tmp992[94], tmp992[93], tmp992[92], tmp992[91], tmp992[90], tmp992[89], tmp992[88], tmp992[87], tmp992[86], tmp992[85], tmp992[84], tmp992[83], tmp992[82], tmp992[81], tmp992[80], tmp992[79], tmp992[78], tmp992[77], tmp992[76], tmp992[75], tmp992[74], tmp992[73], tmp992[72], tmp992[71], tmp992[70], tmp992[69], tmp992[68], tmp992[67], tmp992[66], tmp992[65], tmp992[64], tmp992[63], tmp992[62], tmp992[61], tmp992[60], tmp992[59], tmp992[58], tmp992[57], tmp992[56], tmp992[55], tmp992[54], tmp992[53], tmp992[52], tmp992[51], tmp992[50], tmp992[49], tmp992[48], tmp992[47], tmp992[46], tmp992[45], tmp992[44], tmp992[43], tmp992[42], tmp992[41], tmp992[40], tmp992[39], tmp992[38], tmp992[37], tmp992[36], tmp992[35], tmp992[34], tmp992[33], tmp992[32], tmp992[31], tmp992[30], tmp992[29], tmp992[28], tmp992[27], tmp992[26], tmp992[25], tmp992[24], tmp992[23], tmp992[22], tmp992[21], tmp992[20], tmp992[19], tmp992[18], tmp992[17], tmp992[16], tmp992[15], tmp992[14], tmp992[13], tmp992[12], tmp992[11], tmp992[10], tmp992[9], tmp992[8], tmp992[7], tmp992[6], tmp992[5], tmp992[4], tmp992[3], tmp992[2], tmp992[1], tmp992[0]};
    assign tmp994 = ~tmp35;
    assign tmp995 = ~tmp36;
    assign tmp996 = tmp994 & tmp995;
    assign tmp997 = tmp996 & tmp57;
    assign tmp998 = ~tmp68;
    assign tmp999 = tmp997 & tmp998;
    assign tmp1000 = ~tmp69;
    assign tmp1001 = tmp999 & tmp1000;
    assign tmp1002 = ~tmp108;
    assign tmp1003 = tmp1001 & tmp1002;
    assign tmp1004 = ~tmp375;
    assign tmp1005 = tmp1003 & tmp1004;
    assign tmp1006 = ~tmp470;
    assign tmp1007 = tmp1005 & tmp1006;
    assign tmp1008 = tmp1007 & tmp939;
    assign tmp1009 = tmp16 == _ver_out_tmp_52;
    assign tmp1010 = {const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0, const_113_0};
    assign tmp1011 = {tmp1010, const_112_0};
    assign tmp1012 = tmp1011 - tmp16;
    assign tmp1013 = {const_115_0, const_115_0};
    assign tmp1014 = {tmp1013, const_114_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp1015 = tmp1009 ? tmp1014 : tmp1012;
    assign tmp1016 = {tmp1015[255], tmp1015[254], tmp1015[253], tmp1015[252], tmp1015[251], tmp1015[250], tmp1015[249], tmp1015[248], tmp1015[247], tmp1015[246], tmp1015[245], tmp1015[244], tmp1015[243], tmp1015[242], tmp1015[241], tmp1015[240], tmp1015[239], tmp1015[238], tmp1015[237], tmp1015[236], tmp1015[235], tmp1015[234], tmp1015[233], tmp1015[232], tmp1015[231], tmp1015[230], tmp1015[229], tmp1015[228], tmp1015[227], tmp1015[226], tmp1015[225], tmp1015[224], tmp1015[223], tmp1015[222], tmp1015[221], tmp1015[220], tmp1015[219], tmp1015[218], tmp1015[217], tmp1015[216], tmp1015[215], tmp1015[214], tmp1015[213], tmp1015[212], tmp1015[211], tmp1015[210], tmp1015[209], tmp1015[208], tmp1015[207], tmp1015[206], tmp1015[205], tmp1015[204], tmp1015[203], tmp1015[202], tmp1015[201], tmp1015[200], tmp1015[199], tmp1015[198], tmp1015[197], tmp1015[196], tmp1015[195], tmp1015[194], tmp1015[193], tmp1015[192], tmp1015[191], tmp1015[190], tmp1015[189], tmp1015[188], tmp1015[187], tmp1015[186], tmp1015[185], tmp1015[184], tmp1015[183], tmp1015[182], tmp1015[181], tmp1015[180], tmp1015[179], tmp1015[178], tmp1015[177], tmp1015[176], tmp1015[175], tmp1015[174], tmp1015[173], tmp1015[172], tmp1015[171], tmp1015[170], tmp1015[169], tmp1015[168], tmp1015[167], tmp1015[166], tmp1015[165], tmp1015[164], tmp1015[163], tmp1015[162], tmp1015[161], tmp1015[160], tmp1015[159], tmp1015[158], tmp1015[157], tmp1015[156], tmp1015[155], tmp1015[154], tmp1015[153], tmp1015[152], tmp1015[151], tmp1015[150], tmp1015[149], tmp1015[148], tmp1015[147], tmp1015[146], tmp1015[145], tmp1015[144], tmp1015[143], tmp1015[142], tmp1015[141], tmp1015[140], tmp1015[139], tmp1015[138], tmp1015[137], tmp1015[136], tmp1015[135], tmp1015[134], tmp1015[133], tmp1015[132], tmp1015[131], tmp1015[130], tmp1015[129], tmp1015[128], tmp1015[127], tmp1015[126], tmp1015[125], tmp1015[124], tmp1015[123], tmp1015[122], tmp1015[121], tmp1015[120], tmp1015[119], tmp1015[118], tmp1015[117], tmp1015[116], tmp1015[115], tmp1015[114], tmp1015[113], tmp1015[112], tmp1015[111], tmp1015[110], tmp1015[109], tmp1015[108], tmp1015[107], tmp1015[106], tmp1015[105], tmp1015[104], tmp1015[103], tmp1015[102], tmp1015[101], tmp1015[100], tmp1015[99], tmp1015[98], tmp1015[97], tmp1015[96], tmp1015[95], tmp1015[94], tmp1015[93], tmp1015[92], tmp1015[91], tmp1015[90], tmp1015[89], tmp1015[88], tmp1015[87], tmp1015[86], tmp1015[85], tmp1015[84], tmp1015[83], tmp1015[82], tmp1015[81], tmp1015[80], tmp1015[79], tmp1015[78], tmp1015[77], tmp1015[76], tmp1015[75], tmp1015[74], tmp1015[73], tmp1015[72], tmp1015[71], tmp1015[70], tmp1015[69], tmp1015[68], tmp1015[67], tmp1015[66], tmp1015[65], tmp1015[64], tmp1015[63], tmp1015[62], tmp1015[61], tmp1015[60], tmp1015[59], tmp1015[58], tmp1015[57], tmp1015[56], tmp1015[55], tmp1015[54], tmp1015[53], tmp1015[52], tmp1015[51], tmp1015[50], tmp1015[49], tmp1015[48], tmp1015[47], tmp1015[46], tmp1015[45], tmp1015[44], tmp1015[43], tmp1015[42], tmp1015[41], tmp1015[40], tmp1015[39], tmp1015[38], tmp1015[37], tmp1015[36], tmp1015[35], tmp1015[34], tmp1015[33], tmp1015[32], tmp1015[31], tmp1015[30], tmp1015[29], tmp1015[28], tmp1015[27], tmp1015[26], tmp1015[25], tmp1015[24], tmp1015[23], tmp1015[22], tmp1015[21], tmp1015[20], tmp1015[19], tmp1015[18], tmp1015[17], tmp1015[16], tmp1015[15], tmp1015[14], tmp1015[13], tmp1015[12], tmp1015[11], tmp1015[10], tmp1015[9], tmp1015[8], tmp1015[7], tmp1015[6], tmp1015[5], tmp1015[4], tmp1015[3], tmp1015[2], tmp1015[1], tmp1015[0]};
    assign tmp1017 = ~tmp35;
    assign tmp1018 = ~tmp36;
    assign tmp1019 = tmp1017 & tmp1018;
    assign tmp1020 = tmp1019 & tmp57;
    assign tmp1021 = ~tmp68;
    assign tmp1022 = tmp1020 & tmp1021;
    assign tmp1023 = ~tmp69;
    assign tmp1024 = tmp1022 & tmp1023;
    assign tmp1025 = ~tmp108;
    assign tmp1026 = tmp1024 & tmp1025;
    assign tmp1027 = ~tmp375;
    assign tmp1028 = tmp1026 & tmp1027;
    assign tmp1029 = ~tmp470;
    assign tmp1030 = tmp1028 & tmp1029;
    assign tmp1031 = tmp1030 & tmp939;
    assign tmp1032 = {const_117_0};
    assign tmp1033 = {tmp1032, const_116_2};
    assign tmp1034 = my_calculator_ctrl == tmp1033;
    assign tmp1035 = ~tmp35;
    assign tmp1036 = ~tmp36;
    assign tmp1037 = tmp1035 & tmp1036;
    assign tmp1038 = ~tmp57;
    assign tmp1039 = tmp1037 & tmp1038;
    assign tmp1040 = tmp1039 & tmp1034;
    assign tmp1041 = ~tmp35;
    assign tmp1042 = ~tmp36;
    assign tmp1043 = tmp1041 & tmp1042;
    assign tmp1044 = ~tmp57;
    assign tmp1045 = tmp1043 & tmp1044;
    assign tmp1046 = tmp1045 & tmp1034;
    assign tmp1047 = {const_120_0, const_120_0, const_120_0};
    assign tmp1048 = {tmp1047, const_119_0};
    assign tmp1049 = my_calculator_in_y == tmp1048;
    assign tmp1050 = my_calculator_in_y == const_121_15;
    assign tmp1051 = ~tmp35;
    assign tmp1052 = ~tmp36;
    assign tmp1053 = tmp1051 & tmp1052;
    assign tmp1054 = ~tmp57;
    assign tmp1055 = tmp1053 & tmp1054;
    assign tmp1056 = tmp1055 & tmp1034;
    assign tmp1057 = ~tmp1049;
    assign tmp1058 = tmp1056 & tmp1057;
    assign tmp1059 = tmp1058 & tmp1050;
    assign tmp1060 = ~tmp35;
    assign tmp1061 = ~tmp36;
    assign tmp1062 = tmp1060 & tmp1061;
    assign tmp1063 = ~tmp57;
    assign tmp1064 = tmp1062 & tmp1063;
    assign tmp1065 = tmp1064 & tmp1034;
    assign tmp1066 = ~tmp1049;
    assign tmp1067 = tmp1065 & tmp1066;
    assign tmp1068 = tmp1067 & tmp1050;
    assign tmp1069 = ~tmp35;
    assign tmp1070 = ~tmp36;
    assign tmp1071 = tmp1069 & tmp1070;
    assign tmp1072 = ~tmp57;
    assign tmp1073 = tmp1071 & tmp1072;
    assign tmp1074 = tmp1073 & tmp1034;
    assign tmp1075 = ~tmp1049;
    assign tmp1076 = tmp1074 & tmp1075;
    assign tmp1077 = tmp1076 & tmp1050;
    assign tmp1078 = ~tmp35;
    assign tmp1079 = ~tmp36;
    assign tmp1080 = tmp1078 & tmp1079;
    assign tmp1081 = ~tmp57;
    assign tmp1082 = tmp1080 & tmp1081;
    assign tmp1083 = tmp1082 & tmp1034;
    assign tmp1084 = ~tmp1049;
    assign tmp1085 = tmp1083 & tmp1084;
    assign tmp1086 = tmp1085 & tmp1050;
    assign tmp1087 = {const_123_0, const_123_0, const_123_0};
    assign tmp1088 = {tmp1087, const_122_1};
    assign tmp1089 = my_calculator_in_y == tmp1088;
    assign tmp1090 = {const_125_0, const_125_0};
    assign tmp1091 = {tmp1090, const_124_2};
    assign tmp1092 = my_calculator_in_y == tmp1091;
    assign tmp1093 = tmp1089 | tmp1092;
    assign tmp1094 = {const_127_0, const_127_0};
    assign tmp1095 = {tmp1094, const_126_3};
    assign tmp1096 = my_calculator_in_y == tmp1095;
    assign tmp1097 = tmp1093 | tmp1096;
    assign tmp1098 = {tmp11[254], tmp11[253], tmp11[252], tmp11[251], tmp11[250], tmp11[249], tmp11[248], tmp11[247], tmp11[246], tmp11[245], tmp11[244], tmp11[243], tmp11[242], tmp11[241], tmp11[240], tmp11[239], tmp11[238], tmp11[237], tmp11[236], tmp11[235], tmp11[234], tmp11[233], tmp11[232], tmp11[231], tmp11[230], tmp11[229], tmp11[228], tmp11[227], tmp11[226], tmp11[225], tmp11[224], tmp11[223], tmp11[222], tmp11[221], tmp11[220], tmp11[219], tmp11[218], tmp11[217], tmp11[216], tmp11[215], tmp11[214], tmp11[213], tmp11[212], tmp11[211], tmp11[210], tmp11[209], tmp11[208], tmp11[207], tmp11[206], tmp11[205], tmp11[204], tmp11[203], tmp11[202], tmp11[201], tmp11[200], tmp11[199], tmp11[198], tmp11[197], tmp11[196], tmp11[195], tmp11[194], tmp11[193], tmp11[192], tmp11[191], tmp11[190], tmp11[189], tmp11[188], tmp11[187], tmp11[186], tmp11[185], tmp11[184], tmp11[183], tmp11[182], tmp11[181], tmp11[180], tmp11[179], tmp11[178], tmp11[177], tmp11[176], tmp11[175], tmp11[174], tmp11[173], tmp11[172], tmp11[171], tmp11[170], tmp11[169], tmp11[168], tmp11[167], tmp11[166], tmp11[165], tmp11[164], tmp11[163], tmp11[162], tmp11[161], tmp11[160], tmp11[159], tmp11[158], tmp11[157], tmp11[156], tmp11[155], tmp11[154], tmp11[153], tmp11[152], tmp11[151], tmp11[150], tmp11[149], tmp11[148], tmp11[147], tmp11[146], tmp11[145], tmp11[144], tmp11[143], tmp11[142], tmp11[141], tmp11[140], tmp11[139], tmp11[138], tmp11[137], tmp11[136], tmp11[135], tmp11[134], tmp11[133], tmp11[132], tmp11[131], tmp11[130], tmp11[129], tmp11[128], tmp11[127], tmp11[126], tmp11[125], tmp11[124], tmp11[123], tmp11[122], tmp11[121], tmp11[120], tmp11[119], tmp11[118], tmp11[117], tmp11[116], tmp11[115], tmp11[114], tmp11[113], tmp11[112], tmp11[111], tmp11[110], tmp11[109], tmp11[108], tmp11[107], tmp11[106], tmp11[105], tmp11[104], tmp11[103], tmp11[102], tmp11[101], tmp11[100], tmp11[99], tmp11[98], tmp11[97], tmp11[96], tmp11[95], tmp11[94], tmp11[93], tmp11[92], tmp11[91], tmp11[90], tmp11[89], tmp11[88], tmp11[87], tmp11[86], tmp11[85], tmp11[84], tmp11[83], tmp11[82], tmp11[81], tmp11[80], tmp11[79], tmp11[78], tmp11[77], tmp11[76], tmp11[75], tmp11[74], tmp11[73], tmp11[72], tmp11[71], tmp11[70], tmp11[69], tmp11[68], tmp11[67], tmp11[66], tmp11[65], tmp11[64], tmp11[63], tmp11[62], tmp11[61], tmp11[60], tmp11[59], tmp11[58], tmp11[57], tmp11[56], tmp11[55], tmp11[54], tmp11[53], tmp11[52], tmp11[51], tmp11[50], tmp11[49], tmp11[48], tmp11[47], tmp11[46], tmp11[45], tmp11[44], tmp11[43], tmp11[42], tmp11[41], tmp11[40], tmp11[39], tmp11[38], tmp11[37], tmp11[36], tmp11[35], tmp11[34], tmp11[33], tmp11[32], tmp11[31], tmp11[30], tmp11[29], tmp11[28], tmp11[27], tmp11[26], tmp11[25], tmp11[24], tmp11[23], tmp11[22], tmp11[21], tmp11[20], tmp11[19], tmp11[18], tmp11[17], tmp11[16], tmp11[15], tmp11[14], tmp11[13], tmp11[12], tmp11[11], tmp11[10], tmp11[9], tmp11[8], tmp11[7], tmp11[6], tmp11[5], tmp11[4], tmp11[3], tmp11[2], tmp11[1], tmp11[0]};
    assign tmp1099 = {tmp1098, const_128_0};
    assign tmp1100 = {const_129_0};
    assign tmp1101 = {tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100, tmp1100};
    assign tmp1102 = {tmp1101, const_129_0};
    assign tmp1103 = {tmp11[255]};
    assign tmp1104 = tmp1102 - tmp11;
    assign tmp1105 = {tmp1104[256]};
    assign tmp1106 = {tmp1102[255]};
    assign tmp1107 = ~tmp1106;
    assign tmp1108 = tmp1105 ^ tmp1107;
    assign tmp1109 = {tmp11[255]};
    assign tmp1110 = ~tmp1109;
    assign tmp1111 = tmp1108 ^ tmp1110;
    assign tmp1112 = {tmp1099[255]};
    assign tmp1113 = {const_130_0};
    assign tmp1114 = {tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113, tmp1113};
    assign tmp1115 = {tmp1114, const_130_0};
    assign tmp1116 = tmp1099 - tmp1115;
    assign tmp1117 = {tmp1116[256]};
    assign tmp1118 = {tmp1099[255]};
    assign tmp1119 = ~tmp1118;
    assign tmp1120 = tmp1117 ^ tmp1119;
    assign tmp1121 = {tmp1115[255]};
    assign tmp1122 = ~tmp1121;
    assign tmp1123 = tmp1120 ^ tmp1122;
    assign tmp1124 = tmp1111 & tmp1123;
    assign tmp1125 = {tmp11[255]};
    assign tmp1126 = {const_131_0};
    assign tmp1127 = {tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126, tmp1126};
    assign tmp1128 = {tmp1127, const_131_0};
    assign tmp1129 = tmp11 - tmp1128;
    assign tmp1130 = {tmp1129[256]};
    assign tmp1131 = {tmp11[255]};
    assign tmp1132 = ~tmp1131;
    assign tmp1133 = tmp1130 ^ tmp1132;
    assign tmp1134 = {tmp1128[255]};
    assign tmp1135 = ~tmp1134;
    assign tmp1136 = tmp1133 ^ tmp1135;
    assign tmp1137 = {const_132_0};
    assign tmp1138 = {tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137, tmp1137};
    assign tmp1139 = {tmp1138, const_132_0};
    assign tmp1140 = {tmp1099[255]};
    assign tmp1141 = tmp1139 - tmp1099;
    assign tmp1142 = {tmp1141[256]};
    assign tmp1143 = {tmp1139[255]};
    assign tmp1144 = ~tmp1143;
    assign tmp1145 = tmp1142 ^ tmp1144;
    assign tmp1146 = {tmp1099[255]};
    assign tmp1147 = ~tmp1146;
    assign tmp1148 = tmp1145 ^ tmp1147;
    assign tmp1149 = tmp1139 == tmp1099;
    assign tmp1150 = tmp1148 | tmp1149;
    assign tmp1151 = tmp1136 & tmp1150;
    assign tmp1152 = tmp1124 ? const_133_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp1099;
    assign tmp1153 = tmp1151 ? _ver_out_tmp_60 : tmp1152;
    assign tmp1154 = ~tmp35;
    assign tmp1155 = ~tmp36;
    assign tmp1156 = tmp1154 & tmp1155;
    assign tmp1157 = ~tmp57;
    assign tmp1158 = tmp1156 & tmp1157;
    assign tmp1159 = tmp1158 & tmp1034;
    assign tmp1160 = ~tmp1049;
    assign tmp1161 = tmp1159 & tmp1160;
    assign tmp1162 = ~tmp1050;
    assign tmp1163 = tmp1161 & tmp1162;
    assign tmp1164 = tmp1163 & tmp1097;
    assign tmp1165 = {tmp13[254], tmp13[253], tmp13[252], tmp13[251], tmp13[250], tmp13[249], tmp13[248], tmp13[247], tmp13[246], tmp13[245], tmp13[244], tmp13[243], tmp13[242], tmp13[241], tmp13[240], tmp13[239], tmp13[238], tmp13[237], tmp13[236], tmp13[235], tmp13[234], tmp13[233], tmp13[232], tmp13[231], tmp13[230], tmp13[229], tmp13[228], tmp13[227], tmp13[226], tmp13[225], tmp13[224], tmp13[223], tmp13[222], tmp13[221], tmp13[220], tmp13[219], tmp13[218], tmp13[217], tmp13[216], tmp13[215], tmp13[214], tmp13[213], tmp13[212], tmp13[211], tmp13[210], tmp13[209], tmp13[208], tmp13[207], tmp13[206], tmp13[205], tmp13[204], tmp13[203], tmp13[202], tmp13[201], tmp13[200], tmp13[199], tmp13[198], tmp13[197], tmp13[196], tmp13[195], tmp13[194], tmp13[193], tmp13[192], tmp13[191], tmp13[190], tmp13[189], tmp13[188], tmp13[187], tmp13[186], tmp13[185], tmp13[184], tmp13[183], tmp13[182], tmp13[181], tmp13[180], tmp13[179], tmp13[178], tmp13[177], tmp13[176], tmp13[175], tmp13[174], tmp13[173], tmp13[172], tmp13[171], tmp13[170], tmp13[169], tmp13[168], tmp13[167], tmp13[166], tmp13[165], tmp13[164], tmp13[163], tmp13[162], tmp13[161], tmp13[160], tmp13[159], tmp13[158], tmp13[157], tmp13[156], tmp13[155], tmp13[154], tmp13[153], tmp13[152], tmp13[151], tmp13[150], tmp13[149], tmp13[148], tmp13[147], tmp13[146], tmp13[145], tmp13[144], tmp13[143], tmp13[142], tmp13[141], tmp13[140], tmp13[139], tmp13[138], tmp13[137], tmp13[136], tmp13[135], tmp13[134], tmp13[133], tmp13[132], tmp13[131], tmp13[130], tmp13[129], tmp13[128], tmp13[127], tmp13[126], tmp13[125], tmp13[124], tmp13[123], tmp13[122], tmp13[121], tmp13[120], tmp13[119], tmp13[118], tmp13[117], tmp13[116], tmp13[115], tmp13[114], tmp13[113], tmp13[112], tmp13[111], tmp13[110], tmp13[109], tmp13[108], tmp13[107], tmp13[106], tmp13[105], tmp13[104], tmp13[103], tmp13[102], tmp13[101], tmp13[100], tmp13[99], tmp13[98], tmp13[97], tmp13[96], tmp13[95], tmp13[94], tmp13[93], tmp13[92], tmp13[91], tmp13[90], tmp13[89], tmp13[88], tmp13[87], tmp13[86], tmp13[85], tmp13[84], tmp13[83], tmp13[82], tmp13[81], tmp13[80], tmp13[79], tmp13[78], tmp13[77], tmp13[76], tmp13[75], tmp13[74], tmp13[73], tmp13[72], tmp13[71], tmp13[70], tmp13[69], tmp13[68], tmp13[67], tmp13[66], tmp13[65], tmp13[64], tmp13[63], tmp13[62], tmp13[61], tmp13[60], tmp13[59], tmp13[58], tmp13[57], tmp13[56], tmp13[55], tmp13[54], tmp13[53], tmp13[52], tmp13[51], tmp13[50], tmp13[49], tmp13[48], tmp13[47], tmp13[46], tmp13[45], tmp13[44], tmp13[43], tmp13[42], tmp13[41], tmp13[40], tmp13[39], tmp13[38], tmp13[37], tmp13[36], tmp13[35], tmp13[34], tmp13[33], tmp13[32], tmp13[31], tmp13[30], tmp13[29], tmp13[28], tmp13[27], tmp13[26], tmp13[25], tmp13[24], tmp13[23], tmp13[22], tmp13[21], tmp13[20], tmp13[19], tmp13[18], tmp13[17], tmp13[16], tmp13[15], tmp13[14], tmp13[13], tmp13[12], tmp13[11], tmp13[10], tmp13[9], tmp13[8], tmp13[7], tmp13[6], tmp13[5], tmp13[4], tmp13[3], tmp13[2], tmp13[1], tmp13[0]};
    assign tmp1166 = {tmp1165, const_135_0};
    assign tmp1167 = {const_136_0};
    assign tmp1168 = {tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167, tmp1167};
    assign tmp1169 = {tmp1168, const_136_0};
    assign tmp1170 = {tmp13[255]};
    assign tmp1171 = tmp1169 - tmp13;
    assign tmp1172 = {tmp1171[256]};
    assign tmp1173 = {tmp1169[255]};
    assign tmp1174 = ~tmp1173;
    assign tmp1175 = tmp1172 ^ tmp1174;
    assign tmp1176 = {tmp13[255]};
    assign tmp1177 = ~tmp1176;
    assign tmp1178 = tmp1175 ^ tmp1177;
    assign tmp1179 = {tmp1166[255]};
    assign tmp1180 = {const_137_0};
    assign tmp1181 = {tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180, tmp1180};
    assign tmp1182 = {tmp1181, const_137_0};
    assign tmp1183 = tmp1166 - tmp1182;
    assign tmp1184 = {tmp1183[256]};
    assign tmp1185 = {tmp1166[255]};
    assign tmp1186 = ~tmp1185;
    assign tmp1187 = tmp1184 ^ tmp1186;
    assign tmp1188 = {tmp1182[255]};
    assign tmp1189 = ~tmp1188;
    assign tmp1190 = tmp1187 ^ tmp1189;
    assign tmp1191 = tmp1178 & tmp1190;
    assign tmp1192 = {tmp13[255]};
    assign tmp1193 = {const_138_0};
    assign tmp1194 = {tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193, tmp1193};
    assign tmp1195 = {tmp1194, const_138_0};
    assign tmp1196 = tmp13 - tmp1195;
    assign tmp1197 = {tmp1196[256]};
    assign tmp1198 = {tmp13[255]};
    assign tmp1199 = ~tmp1198;
    assign tmp1200 = tmp1197 ^ tmp1199;
    assign tmp1201 = {tmp1195[255]};
    assign tmp1202 = ~tmp1201;
    assign tmp1203 = tmp1200 ^ tmp1202;
    assign tmp1204 = {const_139_0};
    assign tmp1205 = {tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204, tmp1204};
    assign tmp1206 = {tmp1205, const_139_0};
    assign tmp1207 = {tmp1166[255]};
    assign tmp1208 = tmp1206 - tmp1166;
    assign tmp1209 = {tmp1208[256]};
    assign tmp1210 = {tmp1206[255]};
    assign tmp1211 = ~tmp1210;
    assign tmp1212 = tmp1209 ^ tmp1211;
    assign tmp1213 = {tmp1166[255]};
    assign tmp1214 = ~tmp1213;
    assign tmp1215 = tmp1212 ^ tmp1214;
    assign tmp1216 = tmp1206 == tmp1166;
    assign tmp1217 = tmp1215 | tmp1216;
    assign tmp1218 = tmp1203 & tmp1217;
    assign tmp1219 = tmp1191 ? const_140_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp1166;
    assign tmp1220 = tmp1218 ? _ver_out_tmp_61 : tmp1219;
    assign tmp1221 = ~tmp35;
    assign tmp1222 = ~tmp36;
    assign tmp1223 = tmp1221 & tmp1222;
    assign tmp1224 = ~tmp57;
    assign tmp1225 = tmp1223 & tmp1224;
    assign tmp1226 = tmp1225 & tmp1034;
    assign tmp1227 = ~tmp1049;
    assign tmp1228 = tmp1226 & tmp1227;
    assign tmp1229 = ~tmp1050;
    assign tmp1230 = tmp1228 & tmp1229;
    assign tmp1231 = tmp1230 & tmp1097;
    assign tmp1232 = {tmp15[254], tmp15[253], tmp15[252], tmp15[251], tmp15[250], tmp15[249], tmp15[248], tmp15[247], tmp15[246], tmp15[245], tmp15[244], tmp15[243], tmp15[242], tmp15[241], tmp15[240], tmp15[239], tmp15[238], tmp15[237], tmp15[236], tmp15[235], tmp15[234], tmp15[233], tmp15[232], tmp15[231], tmp15[230], tmp15[229], tmp15[228], tmp15[227], tmp15[226], tmp15[225], tmp15[224], tmp15[223], tmp15[222], tmp15[221], tmp15[220], tmp15[219], tmp15[218], tmp15[217], tmp15[216], tmp15[215], tmp15[214], tmp15[213], tmp15[212], tmp15[211], tmp15[210], tmp15[209], tmp15[208], tmp15[207], tmp15[206], tmp15[205], tmp15[204], tmp15[203], tmp15[202], tmp15[201], tmp15[200], tmp15[199], tmp15[198], tmp15[197], tmp15[196], tmp15[195], tmp15[194], tmp15[193], tmp15[192], tmp15[191], tmp15[190], tmp15[189], tmp15[188], tmp15[187], tmp15[186], tmp15[185], tmp15[184], tmp15[183], tmp15[182], tmp15[181], tmp15[180], tmp15[179], tmp15[178], tmp15[177], tmp15[176], tmp15[175], tmp15[174], tmp15[173], tmp15[172], tmp15[171], tmp15[170], tmp15[169], tmp15[168], tmp15[167], tmp15[166], tmp15[165], tmp15[164], tmp15[163], tmp15[162], tmp15[161], tmp15[160], tmp15[159], tmp15[158], tmp15[157], tmp15[156], tmp15[155], tmp15[154], tmp15[153], tmp15[152], tmp15[151], tmp15[150], tmp15[149], tmp15[148], tmp15[147], tmp15[146], tmp15[145], tmp15[144], tmp15[143], tmp15[142], tmp15[141], tmp15[140], tmp15[139], tmp15[138], tmp15[137], tmp15[136], tmp15[135], tmp15[134], tmp15[133], tmp15[132], tmp15[131], tmp15[130], tmp15[129], tmp15[128], tmp15[127], tmp15[126], tmp15[125], tmp15[124], tmp15[123], tmp15[122], tmp15[121], tmp15[120], tmp15[119], tmp15[118], tmp15[117], tmp15[116], tmp15[115], tmp15[114], tmp15[113], tmp15[112], tmp15[111], tmp15[110], tmp15[109], tmp15[108], tmp15[107], tmp15[106], tmp15[105], tmp15[104], tmp15[103], tmp15[102], tmp15[101], tmp15[100], tmp15[99], tmp15[98], tmp15[97], tmp15[96], tmp15[95], tmp15[94], tmp15[93], tmp15[92], tmp15[91], tmp15[90], tmp15[89], tmp15[88], tmp15[87], tmp15[86], tmp15[85], tmp15[84], tmp15[83], tmp15[82], tmp15[81], tmp15[80], tmp15[79], tmp15[78], tmp15[77], tmp15[76], tmp15[75], tmp15[74], tmp15[73], tmp15[72], tmp15[71], tmp15[70], tmp15[69], tmp15[68], tmp15[67], tmp15[66], tmp15[65], tmp15[64], tmp15[63], tmp15[62], tmp15[61], tmp15[60], tmp15[59], tmp15[58], tmp15[57], tmp15[56], tmp15[55], tmp15[54], tmp15[53], tmp15[52], tmp15[51], tmp15[50], tmp15[49], tmp15[48], tmp15[47], tmp15[46], tmp15[45], tmp15[44], tmp15[43], tmp15[42], tmp15[41], tmp15[40], tmp15[39], tmp15[38], tmp15[37], tmp15[36], tmp15[35], tmp15[34], tmp15[33], tmp15[32], tmp15[31], tmp15[30], tmp15[29], tmp15[28], tmp15[27], tmp15[26], tmp15[25], tmp15[24], tmp15[23], tmp15[22], tmp15[21], tmp15[20], tmp15[19], tmp15[18], tmp15[17], tmp15[16], tmp15[15], tmp15[14], tmp15[13], tmp15[12], tmp15[11], tmp15[10], tmp15[9], tmp15[8], tmp15[7], tmp15[6], tmp15[5], tmp15[4], tmp15[3], tmp15[2], tmp15[1], tmp15[0]};
    assign tmp1233 = {tmp1232, const_142_0};
    assign tmp1234 = {const_143_0};
    assign tmp1235 = {tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234, tmp1234};
    assign tmp1236 = {tmp1235, const_143_0};
    assign tmp1237 = {tmp15[255]};
    assign tmp1238 = tmp1236 - tmp15;
    assign tmp1239 = {tmp1238[256]};
    assign tmp1240 = {tmp1236[255]};
    assign tmp1241 = ~tmp1240;
    assign tmp1242 = tmp1239 ^ tmp1241;
    assign tmp1243 = {tmp15[255]};
    assign tmp1244 = ~tmp1243;
    assign tmp1245 = tmp1242 ^ tmp1244;
    assign tmp1246 = {tmp1233[255]};
    assign tmp1247 = {const_144_0};
    assign tmp1248 = {tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247, tmp1247};
    assign tmp1249 = {tmp1248, const_144_0};
    assign tmp1250 = tmp1233 - tmp1249;
    assign tmp1251 = {tmp1250[256]};
    assign tmp1252 = {tmp1233[255]};
    assign tmp1253 = ~tmp1252;
    assign tmp1254 = tmp1251 ^ tmp1253;
    assign tmp1255 = {tmp1249[255]};
    assign tmp1256 = ~tmp1255;
    assign tmp1257 = tmp1254 ^ tmp1256;
    assign tmp1258 = tmp1245 & tmp1257;
    assign tmp1259 = {tmp15[255]};
    assign tmp1260 = {const_145_0};
    assign tmp1261 = {tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260, tmp1260};
    assign tmp1262 = {tmp1261, const_145_0};
    assign tmp1263 = tmp15 - tmp1262;
    assign tmp1264 = {tmp1263[256]};
    assign tmp1265 = {tmp15[255]};
    assign tmp1266 = ~tmp1265;
    assign tmp1267 = tmp1264 ^ tmp1266;
    assign tmp1268 = {tmp1262[255]};
    assign tmp1269 = ~tmp1268;
    assign tmp1270 = tmp1267 ^ tmp1269;
    assign tmp1271 = {const_146_0};
    assign tmp1272 = {tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271, tmp1271};
    assign tmp1273 = {tmp1272, const_146_0};
    assign tmp1274 = {tmp1233[255]};
    assign tmp1275 = tmp1273 - tmp1233;
    assign tmp1276 = {tmp1275[256]};
    assign tmp1277 = {tmp1273[255]};
    assign tmp1278 = ~tmp1277;
    assign tmp1279 = tmp1276 ^ tmp1278;
    assign tmp1280 = {tmp1233[255]};
    assign tmp1281 = ~tmp1280;
    assign tmp1282 = tmp1279 ^ tmp1281;
    assign tmp1283 = tmp1273 == tmp1233;
    assign tmp1284 = tmp1282 | tmp1283;
    assign tmp1285 = tmp1270 & tmp1284;
    assign tmp1286 = tmp1258 ? const_147_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp1233;
    assign tmp1287 = tmp1285 ? _ver_out_tmp_62 : tmp1286;
    assign tmp1288 = ~tmp35;
    assign tmp1289 = ~tmp36;
    assign tmp1290 = tmp1288 & tmp1289;
    assign tmp1291 = ~tmp57;
    assign tmp1292 = tmp1290 & tmp1291;
    assign tmp1293 = tmp1292 & tmp1034;
    assign tmp1294 = ~tmp1049;
    assign tmp1295 = tmp1293 & tmp1294;
    assign tmp1296 = ~tmp1050;
    assign tmp1297 = tmp1295 & tmp1296;
    assign tmp1298 = tmp1297 & tmp1097;
    assign tmp1299 = {tmp17[254], tmp17[253], tmp17[252], tmp17[251], tmp17[250], tmp17[249], tmp17[248], tmp17[247], tmp17[246], tmp17[245], tmp17[244], tmp17[243], tmp17[242], tmp17[241], tmp17[240], tmp17[239], tmp17[238], tmp17[237], tmp17[236], tmp17[235], tmp17[234], tmp17[233], tmp17[232], tmp17[231], tmp17[230], tmp17[229], tmp17[228], tmp17[227], tmp17[226], tmp17[225], tmp17[224], tmp17[223], tmp17[222], tmp17[221], tmp17[220], tmp17[219], tmp17[218], tmp17[217], tmp17[216], tmp17[215], tmp17[214], tmp17[213], tmp17[212], tmp17[211], tmp17[210], tmp17[209], tmp17[208], tmp17[207], tmp17[206], tmp17[205], tmp17[204], tmp17[203], tmp17[202], tmp17[201], tmp17[200], tmp17[199], tmp17[198], tmp17[197], tmp17[196], tmp17[195], tmp17[194], tmp17[193], tmp17[192], tmp17[191], tmp17[190], tmp17[189], tmp17[188], tmp17[187], tmp17[186], tmp17[185], tmp17[184], tmp17[183], tmp17[182], tmp17[181], tmp17[180], tmp17[179], tmp17[178], tmp17[177], tmp17[176], tmp17[175], tmp17[174], tmp17[173], tmp17[172], tmp17[171], tmp17[170], tmp17[169], tmp17[168], tmp17[167], tmp17[166], tmp17[165], tmp17[164], tmp17[163], tmp17[162], tmp17[161], tmp17[160], tmp17[159], tmp17[158], tmp17[157], tmp17[156], tmp17[155], tmp17[154], tmp17[153], tmp17[152], tmp17[151], tmp17[150], tmp17[149], tmp17[148], tmp17[147], tmp17[146], tmp17[145], tmp17[144], tmp17[143], tmp17[142], tmp17[141], tmp17[140], tmp17[139], tmp17[138], tmp17[137], tmp17[136], tmp17[135], tmp17[134], tmp17[133], tmp17[132], tmp17[131], tmp17[130], tmp17[129], tmp17[128], tmp17[127], tmp17[126], tmp17[125], tmp17[124], tmp17[123], tmp17[122], tmp17[121], tmp17[120], tmp17[119], tmp17[118], tmp17[117], tmp17[116], tmp17[115], tmp17[114], tmp17[113], tmp17[112], tmp17[111], tmp17[110], tmp17[109], tmp17[108], tmp17[107], tmp17[106], tmp17[105], tmp17[104], tmp17[103], tmp17[102], tmp17[101], tmp17[100], tmp17[99], tmp17[98], tmp17[97], tmp17[96], tmp17[95], tmp17[94], tmp17[93], tmp17[92], tmp17[91], tmp17[90], tmp17[89], tmp17[88], tmp17[87], tmp17[86], tmp17[85], tmp17[84], tmp17[83], tmp17[82], tmp17[81], tmp17[80], tmp17[79], tmp17[78], tmp17[77], tmp17[76], tmp17[75], tmp17[74], tmp17[73], tmp17[72], tmp17[71], tmp17[70], tmp17[69], tmp17[68], tmp17[67], tmp17[66], tmp17[65], tmp17[64], tmp17[63], tmp17[62], tmp17[61], tmp17[60], tmp17[59], tmp17[58], tmp17[57], tmp17[56], tmp17[55], tmp17[54], tmp17[53], tmp17[52], tmp17[51], tmp17[50], tmp17[49], tmp17[48], tmp17[47], tmp17[46], tmp17[45], tmp17[44], tmp17[43], tmp17[42], tmp17[41], tmp17[40], tmp17[39], tmp17[38], tmp17[37], tmp17[36], tmp17[35], tmp17[34], tmp17[33], tmp17[32], tmp17[31], tmp17[30], tmp17[29], tmp17[28], tmp17[27], tmp17[26], tmp17[25], tmp17[24], tmp17[23], tmp17[22], tmp17[21], tmp17[20], tmp17[19], tmp17[18], tmp17[17], tmp17[16], tmp17[15], tmp17[14], tmp17[13], tmp17[12], tmp17[11], tmp17[10], tmp17[9], tmp17[8], tmp17[7], tmp17[6], tmp17[5], tmp17[4], tmp17[3], tmp17[2], tmp17[1], tmp17[0]};
    assign tmp1300 = {tmp1299, const_149_0};
    assign tmp1301 = {const_150_0};
    assign tmp1302 = {tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301, tmp1301};
    assign tmp1303 = {tmp1302, const_150_0};
    assign tmp1304 = {tmp17[255]};
    assign tmp1305 = tmp1303 - tmp17;
    assign tmp1306 = {tmp1305[256]};
    assign tmp1307 = {tmp1303[255]};
    assign tmp1308 = ~tmp1307;
    assign tmp1309 = tmp1306 ^ tmp1308;
    assign tmp1310 = {tmp17[255]};
    assign tmp1311 = ~tmp1310;
    assign tmp1312 = tmp1309 ^ tmp1311;
    assign tmp1313 = {tmp1300[255]};
    assign tmp1314 = {const_151_0};
    assign tmp1315 = {tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314, tmp1314};
    assign tmp1316 = {tmp1315, const_151_0};
    assign tmp1317 = tmp1300 - tmp1316;
    assign tmp1318 = {tmp1317[256]};
    assign tmp1319 = {tmp1300[255]};
    assign tmp1320 = ~tmp1319;
    assign tmp1321 = tmp1318 ^ tmp1320;
    assign tmp1322 = {tmp1316[255]};
    assign tmp1323 = ~tmp1322;
    assign tmp1324 = tmp1321 ^ tmp1323;
    assign tmp1325 = tmp1312 & tmp1324;
    assign tmp1326 = {tmp17[255]};
    assign tmp1327 = {const_152_0};
    assign tmp1328 = {tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327, tmp1327};
    assign tmp1329 = {tmp1328, const_152_0};
    assign tmp1330 = tmp17 - tmp1329;
    assign tmp1331 = {tmp1330[256]};
    assign tmp1332 = {tmp17[255]};
    assign tmp1333 = ~tmp1332;
    assign tmp1334 = tmp1331 ^ tmp1333;
    assign tmp1335 = {tmp1329[255]};
    assign tmp1336 = ~tmp1335;
    assign tmp1337 = tmp1334 ^ tmp1336;
    assign tmp1338 = {const_153_0};
    assign tmp1339 = {tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338, tmp1338};
    assign tmp1340 = {tmp1339, const_153_0};
    assign tmp1341 = {tmp1300[255]};
    assign tmp1342 = tmp1340 - tmp1300;
    assign tmp1343 = {tmp1342[256]};
    assign tmp1344 = {tmp1340[255]};
    assign tmp1345 = ~tmp1344;
    assign tmp1346 = tmp1343 ^ tmp1345;
    assign tmp1347 = {tmp1300[255]};
    assign tmp1348 = ~tmp1347;
    assign tmp1349 = tmp1346 ^ tmp1348;
    assign tmp1350 = tmp1340 == tmp1300;
    assign tmp1351 = tmp1349 | tmp1350;
    assign tmp1352 = tmp1337 & tmp1351;
    assign tmp1353 = tmp1325 ? const_154_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp1300;
    assign tmp1354 = tmp1352 ? _ver_out_tmp_64 : tmp1353;
    assign tmp1355 = ~tmp35;
    assign tmp1356 = ~tmp36;
    assign tmp1357 = tmp1355 & tmp1356;
    assign tmp1358 = ~tmp57;
    assign tmp1359 = tmp1357 & tmp1358;
    assign tmp1360 = tmp1359 & tmp1034;
    assign tmp1361 = ~tmp1049;
    assign tmp1362 = tmp1360 & tmp1361;
    assign tmp1363 = ~tmp1050;
    assign tmp1364 = tmp1362 & tmp1363;
    assign tmp1365 = tmp1364 & tmp1097;
    assign tmp1366 = {const_157_0};
    assign tmp1367 = {tmp1366, const_156_6};
    assign tmp1368 = my_calculator_in_y == tmp1367;
    assign tmp1369 = {const_159_0};
    assign tmp1370 = {tmp1369, const_158_7};
    assign tmp1371 = my_calculator_in_y == tmp1370;
    assign tmp1372 = tmp1368 | tmp1371;
    assign tmp1373 = ~tmp35;
    assign tmp1374 = ~tmp36;
    assign tmp1375 = tmp1373 & tmp1374;
    assign tmp1376 = ~tmp57;
    assign tmp1377 = tmp1375 & tmp1376;
    assign tmp1378 = tmp1377 & tmp1034;
    assign tmp1379 = ~tmp1049;
    assign tmp1380 = tmp1378 & tmp1379;
    assign tmp1381 = ~tmp1050;
    assign tmp1382 = tmp1380 & tmp1381;
    assign tmp1383 = ~tmp1097;
    assign tmp1384 = tmp1382 & tmp1383;
    assign tmp1385 = tmp1384 & tmp1372;
    assign tmp1386 = ~tmp35;
    assign tmp1387 = ~tmp36;
    assign tmp1388 = tmp1386 & tmp1387;
    assign tmp1389 = ~tmp57;
    assign tmp1390 = tmp1388 & tmp1389;
    assign tmp1391 = tmp1390 & tmp1034;
    assign tmp1392 = ~tmp1049;
    assign tmp1393 = tmp1391 & tmp1392;
    assign tmp1394 = ~tmp1050;
    assign tmp1395 = tmp1393 & tmp1394;
    assign tmp1396 = ~tmp1097;
    assign tmp1397 = tmp1395 & tmp1396;
    assign tmp1398 = tmp1397 & tmp1372;
    assign tmp1399 = ~tmp35;
    assign tmp1400 = ~tmp36;
    assign tmp1401 = tmp1399 & tmp1400;
    assign tmp1402 = ~tmp57;
    assign tmp1403 = tmp1401 & tmp1402;
    assign tmp1404 = tmp1403 & tmp1034;
    assign tmp1405 = ~tmp1049;
    assign tmp1406 = tmp1404 & tmp1405;
    assign tmp1407 = ~tmp1050;
    assign tmp1408 = tmp1406 & tmp1407;
    assign tmp1409 = ~tmp1097;
    assign tmp1410 = tmp1408 & tmp1409;
    assign tmp1411 = tmp1410 & tmp1372;
    assign tmp1412 = ~tmp35;
    assign tmp1413 = ~tmp36;
    assign tmp1414 = tmp1412 & tmp1413;
    assign tmp1415 = ~tmp57;
    assign tmp1416 = tmp1414 & tmp1415;
    assign tmp1417 = tmp1416 & tmp1034;
    assign tmp1418 = ~tmp1049;
    assign tmp1419 = tmp1417 & tmp1418;
    assign tmp1420 = ~tmp1050;
    assign tmp1421 = tmp1419 & tmp1420;
    assign tmp1422 = ~tmp1097;
    assign tmp1423 = tmp1421 & tmp1422;
    assign tmp1424 = tmp1423 & tmp1372;
    assign tmp1425 = ~tmp35;
    assign tmp1426 = ~tmp36;
    assign tmp1427 = tmp1425 & tmp1426;
    assign tmp1428 = ~tmp57;
    assign tmp1429 = tmp1427 & tmp1428;
    assign tmp1430 = tmp1429 & tmp1034;
    assign tmp1431 = ~tmp1049;
    assign tmp1432 = tmp1430 & tmp1431;
    assign tmp1433 = ~tmp1050;
    assign tmp1434 = tmp1432 & tmp1433;
    assign tmp1435 = ~tmp1097;
    assign tmp1436 = tmp1434 & tmp1435;
    assign tmp1437 = tmp1436 & tmp1372;
    assign tmp1438 = ~tmp35;
    assign tmp1439 = ~tmp36;
    assign tmp1440 = tmp1438 & tmp1439;
    assign tmp1441 = ~tmp57;
    assign tmp1442 = tmp1440 & tmp1441;
    assign tmp1443 = tmp1442 & tmp1034;
    assign tmp1444 = ~tmp1049;
    assign tmp1445 = tmp1443 & tmp1444;
    assign tmp1446 = ~tmp1050;
    assign tmp1447 = tmp1445 & tmp1446;
    assign tmp1448 = ~tmp1097;
    assign tmp1449 = tmp1447 & tmp1448;
    assign tmp1450 = tmp1449 & tmp1372;
    assign tmp1451 = ~tmp35;
    assign tmp1452 = ~tmp36;
    assign tmp1453 = tmp1451 & tmp1452;
    assign tmp1454 = ~tmp57;
    assign tmp1455 = tmp1453 & tmp1454;
    assign tmp1456 = tmp1455 & tmp1034;
    assign tmp1457 = ~tmp1049;
    assign tmp1458 = tmp1456 & tmp1457;
    assign tmp1459 = ~tmp1050;
    assign tmp1460 = tmp1458 & tmp1459;
    assign tmp1461 = ~tmp1097;
    assign tmp1462 = tmp1460 & tmp1461;
    assign tmp1463 = tmp1462 & tmp1372;
    assign tmp1464 = ~tmp35;
    assign tmp1465 = ~tmp36;
    assign tmp1466 = tmp1464 & tmp1465;
    assign tmp1467 = ~tmp57;
    assign tmp1468 = tmp1466 & tmp1467;
    assign tmp1469 = tmp1468 & tmp1034;
    assign tmp1470 = ~tmp1049;
    assign tmp1471 = tmp1469 & tmp1470;
    assign tmp1472 = ~tmp1050;
    assign tmp1473 = tmp1471 & tmp1472;
    assign tmp1474 = ~tmp1097;
    assign tmp1475 = tmp1473 & tmp1474;
    assign tmp1476 = tmp1475 & tmp1372;
    assign tmp1477 = {const_161_0};
    assign tmp1478 = {tmp1477, const_160_4};
    assign tmp1479 = my_calculator_in_y == tmp1478;
    assign tmp1480 = {const_163_0};
    assign tmp1481 = {tmp1480, const_162_5};
    assign tmp1482 = my_calculator_in_y == tmp1481;
    assign tmp1483 = tmp1479 | tmp1482;
    assign tmp1484 = {tmp11[255]};
    assign tmp1485 = {tmp1484};
    assign tmp1486 = {tmp1485, tmp11};
    assign tmp1487 = {tmp12[255]};
    assign tmp1488 = {tmp1487};
    assign tmp1489 = {tmp1488, tmp12};
    assign tmp1490 = tmp1486 + tmp1489;
    assign tmp1491 = {tmp1490[256], tmp1490[255], tmp1490[254], tmp1490[253], tmp1490[252], tmp1490[251], tmp1490[250], tmp1490[249], tmp1490[248], tmp1490[247], tmp1490[246], tmp1490[245], tmp1490[244], tmp1490[243], tmp1490[242], tmp1490[241], tmp1490[240], tmp1490[239], tmp1490[238], tmp1490[237], tmp1490[236], tmp1490[235], tmp1490[234], tmp1490[233], tmp1490[232], tmp1490[231], tmp1490[230], tmp1490[229], tmp1490[228], tmp1490[227], tmp1490[226], tmp1490[225], tmp1490[224], tmp1490[223], tmp1490[222], tmp1490[221], tmp1490[220], tmp1490[219], tmp1490[218], tmp1490[217], tmp1490[216], tmp1490[215], tmp1490[214], tmp1490[213], tmp1490[212], tmp1490[211], tmp1490[210], tmp1490[209], tmp1490[208], tmp1490[207], tmp1490[206], tmp1490[205], tmp1490[204], tmp1490[203], tmp1490[202], tmp1490[201], tmp1490[200], tmp1490[199], tmp1490[198], tmp1490[197], tmp1490[196], tmp1490[195], tmp1490[194], tmp1490[193], tmp1490[192], tmp1490[191], tmp1490[190], tmp1490[189], tmp1490[188], tmp1490[187], tmp1490[186], tmp1490[185], tmp1490[184], tmp1490[183], tmp1490[182], tmp1490[181], tmp1490[180], tmp1490[179], tmp1490[178], tmp1490[177], tmp1490[176], tmp1490[175], tmp1490[174], tmp1490[173], tmp1490[172], tmp1490[171], tmp1490[170], tmp1490[169], tmp1490[168], tmp1490[167], tmp1490[166], tmp1490[165], tmp1490[164], tmp1490[163], tmp1490[162], tmp1490[161], tmp1490[160], tmp1490[159], tmp1490[158], tmp1490[157], tmp1490[156], tmp1490[155], tmp1490[154], tmp1490[153], tmp1490[152], tmp1490[151], tmp1490[150], tmp1490[149], tmp1490[148], tmp1490[147], tmp1490[146], tmp1490[145], tmp1490[144], tmp1490[143], tmp1490[142], tmp1490[141], tmp1490[140], tmp1490[139], tmp1490[138], tmp1490[137], tmp1490[136], tmp1490[135], tmp1490[134], tmp1490[133], tmp1490[132], tmp1490[131], tmp1490[130], tmp1490[129], tmp1490[128], tmp1490[127], tmp1490[126], tmp1490[125], tmp1490[124], tmp1490[123], tmp1490[122], tmp1490[121], tmp1490[120], tmp1490[119], tmp1490[118], tmp1490[117], tmp1490[116], tmp1490[115], tmp1490[114], tmp1490[113], tmp1490[112], tmp1490[111], tmp1490[110], tmp1490[109], tmp1490[108], tmp1490[107], tmp1490[106], tmp1490[105], tmp1490[104], tmp1490[103], tmp1490[102], tmp1490[101], tmp1490[100], tmp1490[99], tmp1490[98], tmp1490[97], tmp1490[96], tmp1490[95], tmp1490[94], tmp1490[93], tmp1490[92], tmp1490[91], tmp1490[90], tmp1490[89], tmp1490[88], tmp1490[87], tmp1490[86], tmp1490[85], tmp1490[84], tmp1490[83], tmp1490[82], tmp1490[81], tmp1490[80], tmp1490[79], tmp1490[78], tmp1490[77], tmp1490[76], tmp1490[75], tmp1490[74], tmp1490[73], tmp1490[72], tmp1490[71], tmp1490[70], tmp1490[69], tmp1490[68], tmp1490[67], tmp1490[66], tmp1490[65], tmp1490[64], tmp1490[63], tmp1490[62], tmp1490[61], tmp1490[60], tmp1490[59], tmp1490[58], tmp1490[57], tmp1490[56], tmp1490[55], tmp1490[54], tmp1490[53], tmp1490[52], tmp1490[51], tmp1490[50], tmp1490[49], tmp1490[48], tmp1490[47], tmp1490[46], tmp1490[45], tmp1490[44], tmp1490[43], tmp1490[42], tmp1490[41], tmp1490[40], tmp1490[39], tmp1490[38], tmp1490[37], tmp1490[36], tmp1490[35], tmp1490[34], tmp1490[33], tmp1490[32], tmp1490[31], tmp1490[30], tmp1490[29], tmp1490[28], tmp1490[27], tmp1490[26], tmp1490[25], tmp1490[24], tmp1490[23], tmp1490[22], tmp1490[21], tmp1490[20], tmp1490[19], tmp1490[18], tmp1490[17], tmp1490[16], tmp1490[15], tmp1490[14], tmp1490[13], tmp1490[12], tmp1490[11], tmp1490[10], tmp1490[9], tmp1490[8], tmp1490[7], tmp1490[6], tmp1490[5], tmp1490[4], tmp1490[3], tmp1490[2], tmp1490[1], tmp1490[0]};
    assign tmp1492 = {tmp1491[255], tmp1491[254], tmp1491[253], tmp1491[252], tmp1491[251], tmp1491[250], tmp1491[249], tmp1491[248], tmp1491[247], tmp1491[246], tmp1491[245], tmp1491[244], tmp1491[243], tmp1491[242], tmp1491[241], tmp1491[240], tmp1491[239], tmp1491[238], tmp1491[237], tmp1491[236], tmp1491[235], tmp1491[234], tmp1491[233], tmp1491[232], tmp1491[231], tmp1491[230], tmp1491[229], tmp1491[228], tmp1491[227], tmp1491[226], tmp1491[225], tmp1491[224], tmp1491[223], tmp1491[222], tmp1491[221], tmp1491[220], tmp1491[219], tmp1491[218], tmp1491[217], tmp1491[216], tmp1491[215], tmp1491[214], tmp1491[213], tmp1491[212], tmp1491[211], tmp1491[210], tmp1491[209], tmp1491[208], tmp1491[207], tmp1491[206], tmp1491[205], tmp1491[204], tmp1491[203], tmp1491[202], tmp1491[201], tmp1491[200], tmp1491[199], tmp1491[198], tmp1491[197], tmp1491[196], tmp1491[195], tmp1491[194], tmp1491[193], tmp1491[192], tmp1491[191], tmp1491[190], tmp1491[189], tmp1491[188], tmp1491[187], tmp1491[186], tmp1491[185], tmp1491[184], tmp1491[183], tmp1491[182], tmp1491[181], tmp1491[180], tmp1491[179], tmp1491[178], tmp1491[177], tmp1491[176], tmp1491[175], tmp1491[174], tmp1491[173], tmp1491[172], tmp1491[171], tmp1491[170], tmp1491[169], tmp1491[168], tmp1491[167], tmp1491[166], tmp1491[165], tmp1491[164], tmp1491[163], tmp1491[162], tmp1491[161], tmp1491[160], tmp1491[159], tmp1491[158], tmp1491[157], tmp1491[156], tmp1491[155], tmp1491[154], tmp1491[153], tmp1491[152], tmp1491[151], tmp1491[150], tmp1491[149], tmp1491[148], tmp1491[147], tmp1491[146], tmp1491[145], tmp1491[144], tmp1491[143], tmp1491[142], tmp1491[141], tmp1491[140], tmp1491[139], tmp1491[138], tmp1491[137], tmp1491[136], tmp1491[135], tmp1491[134], tmp1491[133], tmp1491[132], tmp1491[131], tmp1491[130], tmp1491[129], tmp1491[128], tmp1491[127], tmp1491[126], tmp1491[125], tmp1491[124], tmp1491[123], tmp1491[122], tmp1491[121], tmp1491[120], tmp1491[119], tmp1491[118], tmp1491[117], tmp1491[116], tmp1491[115], tmp1491[114], tmp1491[113], tmp1491[112], tmp1491[111], tmp1491[110], tmp1491[109], tmp1491[108], tmp1491[107], tmp1491[106], tmp1491[105], tmp1491[104], tmp1491[103], tmp1491[102], tmp1491[101], tmp1491[100], tmp1491[99], tmp1491[98], tmp1491[97], tmp1491[96], tmp1491[95], tmp1491[94], tmp1491[93], tmp1491[92], tmp1491[91], tmp1491[90], tmp1491[89], tmp1491[88], tmp1491[87], tmp1491[86], tmp1491[85], tmp1491[84], tmp1491[83], tmp1491[82], tmp1491[81], tmp1491[80], tmp1491[79], tmp1491[78], tmp1491[77], tmp1491[76], tmp1491[75], tmp1491[74], tmp1491[73], tmp1491[72], tmp1491[71], tmp1491[70], tmp1491[69], tmp1491[68], tmp1491[67], tmp1491[66], tmp1491[65], tmp1491[64], tmp1491[63], tmp1491[62], tmp1491[61], tmp1491[60], tmp1491[59], tmp1491[58], tmp1491[57], tmp1491[56], tmp1491[55], tmp1491[54], tmp1491[53], tmp1491[52], tmp1491[51], tmp1491[50], tmp1491[49], tmp1491[48], tmp1491[47], tmp1491[46], tmp1491[45], tmp1491[44], tmp1491[43], tmp1491[42], tmp1491[41], tmp1491[40], tmp1491[39], tmp1491[38], tmp1491[37], tmp1491[36], tmp1491[35], tmp1491[34], tmp1491[33], tmp1491[32], tmp1491[31], tmp1491[30], tmp1491[29], tmp1491[28], tmp1491[27], tmp1491[26], tmp1491[25], tmp1491[24], tmp1491[23], tmp1491[22], tmp1491[21], tmp1491[20], tmp1491[19], tmp1491[18], tmp1491[17], tmp1491[16], tmp1491[15], tmp1491[14], tmp1491[13], tmp1491[12], tmp1491[11], tmp1491[10], tmp1491[9], tmp1491[8], tmp1491[7], tmp1491[6], tmp1491[5], tmp1491[4], tmp1491[3], tmp1491[2], tmp1491[1], tmp1491[0]};
    assign tmp1493 = {const_164_0};
    assign tmp1494 = {tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493, tmp1493};
    assign tmp1495 = {tmp1494, const_164_0};
    assign tmp1496 = {tmp11[255]};
    assign tmp1497 = tmp1495 - tmp11;
    assign tmp1498 = {tmp1497[256]};
    assign tmp1499 = {tmp1495[255]};
    assign tmp1500 = ~tmp1499;
    assign tmp1501 = tmp1498 ^ tmp1500;
    assign tmp1502 = {tmp11[255]};
    assign tmp1503 = ~tmp1502;
    assign tmp1504 = tmp1501 ^ tmp1503;
    assign tmp1505 = {const_165_0};
    assign tmp1506 = {tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505, tmp1505};
    assign tmp1507 = {tmp1506, const_165_0};
    assign tmp1508 = {tmp12[255]};
    assign tmp1509 = tmp1507 - tmp12;
    assign tmp1510 = {tmp1509[256]};
    assign tmp1511 = {tmp1507[255]};
    assign tmp1512 = ~tmp1511;
    assign tmp1513 = tmp1510 ^ tmp1512;
    assign tmp1514 = {tmp12[255]};
    assign tmp1515 = ~tmp1514;
    assign tmp1516 = tmp1513 ^ tmp1515;
    assign tmp1517 = tmp1504 & tmp1516;
    assign tmp1518 = {tmp1492[255]};
    assign tmp1519 = {const_166_0};
    assign tmp1520 = {tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519, tmp1519};
    assign tmp1521 = {tmp1520, const_166_0};
    assign tmp1522 = tmp1492 - tmp1521;
    assign tmp1523 = {tmp1522[256]};
    assign tmp1524 = {tmp1492[255]};
    assign tmp1525 = ~tmp1524;
    assign tmp1526 = tmp1523 ^ tmp1525;
    assign tmp1527 = {tmp1521[255]};
    assign tmp1528 = ~tmp1527;
    assign tmp1529 = tmp1526 ^ tmp1528;
    assign tmp1530 = tmp1492 == tmp1521;
    assign tmp1531 = tmp1529 | tmp1530;
    assign tmp1532 = tmp1517 & tmp1531;
    assign tmp1533 = {tmp11[255]};
    assign tmp1534 = {const_167_0};
    assign tmp1535 = {tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534, tmp1534};
    assign tmp1536 = {tmp1535, const_167_0};
    assign tmp1537 = tmp11 - tmp1536;
    assign tmp1538 = {tmp1537[256]};
    assign tmp1539 = {tmp11[255]};
    assign tmp1540 = ~tmp1539;
    assign tmp1541 = tmp1538 ^ tmp1540;
    assign tmp1542 = {tmp1536[255]};
    assign tmp1543 = ~tmp1542;
    assign tmp1544 = tmp1541 ^ tmp1543;
    assign tmp1545 = {tmp12[255]};
    assign tmp1546 = {const_168_0};
    assign tmp1547 = {tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546, tmp1546};
    assign tmp1548 = {tmp1547, const_168_0};
    assign tmp1549 = tmp12 - tmp1548;
    assign tmp1550 = {tmp1549[256]};
    assign tmp1551 = {tmp12[255]};
    assign tmp1552 = ~tmp1551;
    assign tmp1553 = tmp1550 ^ tmp1552;
    assign tmp1554 = {tmp1548[255]};
    assign tmp1555 = ~tmp1554;
    assign tmp1556 = tmp1553 ^ tmp1555;
    assign tmp1557 = tmp1544 & tmp1556;
    assign tmp1558 = {const_169_0};
    assign tmp1559 = {tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558, tmp1558};
    assign tmp1560 = {tmp1559, const_169_0};
    assign tmp1561 = {tmp1492[255]};
    assign tmp1562 = tmp1560 - tmp1492;
    assign tmp1563 = {tmp1562[256]};
    assign tmp1564 = {tmp1560[255]};
    assign tmp1565 = ~tmp1564;
    assign tmp1566 = tmp1563 ^ tmp1565;
    assign tmp1567 = {tmp1492[255]};
    assign tmp1568 = ~tmp1567;
    assign tmp1569 = tmp1566 ^ tmp1568;
    assign tmp1570 = tmp1560 == tmp1492;
    assign tmp1571 = tmp1569 | tmp1570;
    assign tmp1572 = tmp1557 & tmp1571;
    assign tmp1573 = tmp1532 ? const_170_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp1492;
    assign tmp1574 = tmp1572 ? _ver_out_tmp_67 : tmp1573;
    assign tmp1575 = ~tmp35;
    assign tmp1576 = ~tmp36;
    assign tmp1577 = tmp1575 & tmp1576;
    assign tmp1578 = ~tmp57;
    assign tmp1579 = tmp1577 & tmp1578;
    assign tmp1580 = tmp1579 & tmp1034;
    assign tmp1581 = ~tmp1049;
    assign tmp1582 = tmp1580 & tmp1581;
    assign tmp1583 = ~tmp1050;
    assign tmp1584 = tmp1582 & tmp1583;
    assign tmp1585 = ~tmp1097;
    assign tmp1586 = tmp1584 & tmp1585;
    assign tmp1587 = ~tmp1372;
    assign tmp1588 = tmp1586 & tmp1587;
    assign tmp1589 = tmp1588 & tmp1483;
    assign tmp1590 = ~tmp35;
    assign tmp1591 = ~tmp36;
    assign tmp1592 = tmp1590 & tmp1591;
    assign tmp1593 = ~tmp57;
    assign tmp1594 = tmp1592 & tmp1593;
    assign tmp1595 = tmp1594 & tmp1034;
    assign tmp1596 = ~tmp1049;
    assign tmp1597 = tmp1595 & tmp1596;
    assign tmp1598 = ~tmp1050;
    assign tmp1599 = tmp1597 & tmp1598;
    assign tmp1600 = ~tmp1097;
    assign tmp1601 = tmp1599 & tmp1600;
    assign tmp1602 = ~tmp1372;
    assign tmp1603 = tmp1601 & tmp1602;
    assign tmp1604 = tmp1603 & tmp1483;
    assign tmp1605 = {tmp13[255]};
    assign tmp1606 = {tmp1605};
    assign tmp1607 = {tmp1606, tmp13};
    assign tmp1608 = {tmp14[255]};
    assign tmp1609 = {tmp1608};
    assign tmp1610 = {tmp1609, tmp14};
    assign tmp1611 = tmp1607 + tmp1610;
    assign tmp1612 = {tmp1611[256], tmp1611[255], tmp1611[254], tmp1611[253], tmp1611[252], tmp1611[251], tmp1611[250], tmp1611[249], tmp1611[248], tmp1611[247], tmp1611[246], tmp1611[245], tmp1611[244], tmp1611[243], tmp1611[242], tmp1611[241], tmp1611[240], tmp1611[239], tmp1611[238], tmp1611[237], tmp1611[236], tmp1611[235], tmp1611[234], tmp1611[233], tmp1611[232], tmp1611[231], tmp1611[230], tmp1611[229], tmp1611[228], tmp1611[227], tmp1611[226], tmp1611[225], tmp1611[224], tmp1611[223], tmp1611[222], tmp1611[221], tmp1611[220], tmp1611[219], tmp1611[218], tmp1611[217], tmp1611[216], tmp1611[215], tmp1611[214], tmp1611[213], tmp1611[212], tmp1611[211], tmp1611[210], tmp1611[209], tmp1611[208], tmp1611[207], tmp1611[206], tmp1611[205], tmp1611[204], tmp1611[203], tmp1611[202], tmp1611[201], tmp1611[200], tmp1611[199], tmp1611[198], tmp1611[197], tmp1611[196], tmp1611[195], tmp1611[194], tmp1611[193], tmp1611[192], tmp1611[191], tmp1611[190], tmp1611[189], tmp1611[188], tmp1611[187], tmp1611[186], tmp1611[185], tmp1611[184], tmp1611[183], tmp1611[182], tmp1611[181], tmp1611[180], tmp1611[179], tmp1611[178], tmp1611[177], tmp1611[176], tmp1611[175], tmp1611[174], tmp1611[173], tmp1611[172], tmp1611[171], tmp1611[170], tmp1611[169], tmp1611[168], tmp1611[167], tmp1611[166], tmp1611[165], tmp1611[164], tmp1611[163], tmp1611[162], tmp1611[161], tmp1611[160], tmp1611[159], tmp1611[158], tmp1611[157], tmp1611[156], tmp1611[155], tmp1611[154], tmp1611[153], tmp1611[152], tmp1611[151], tmp1611[150], tmp1611[149], tmp1611[148], tmp1611[147], tmp1611[146], tmp1611[145], tmp1611[144], tmp1611[143], tmp1611[142], tmp1611[141], tmp1611[140], tmp1611[139], tmp1611[138], tmp1611[137], tmp1611[136], tmp1611[135], tmp1611[134], tmp1611[133], tmp1611[132], tmp1611[131], tmp1611[130], tmp1611[129], tmp1611[128], tmp1611[127], tmp1611[126], tmp1611[125], tmp1611[124], tmp1611[123], tmp1611[122], tmp1611[121], tmp1611[120], tmp1611[119], tmp1611[118], tmp1611[117], tmp1611[116], tmp1611[115], tmp1611[114], tmp1611[113], tmp1611[112], tmp1611[111], tmp1611[110], tmp1611[109], tmp1611[108], tmp1611[107], tmp1611[106], tmp1611[105], tmp1611[104], tmp1611[103], tmp1611[102], tmp1611[101], tmp1611[100], tmp1611[99], tmp1611[98], tmp1611[97], tmp1611[96], tmp1611[95], tmp1611[94], tmp1611[93], tmp1611[92], tmp1611[91], tmp1611[90], tmp1611[89], tmp1611[88], tmp1611[87], tmp1611[86], tmp1611[85], tmp1611[84], tmp1611[83], tmp1611[82], tmp1611[81], tmp1611[80], tmp1611[79], tmp1611[78], tmp1611[77], tmp1611[76], tmp1611[75], tmp1611[74], tmp1611[73], tmp1611[72], tmp1611[71], tmp1611[70], tmp1611[69], tmp1611[68], tmp1611[67], tmp1611[66], tmp1611[65], tmp1611[64], tmp1611[63], tmp1611[62], tmp1611[61], tmp1611[60], tmp1611[59], tmp1611[58], tmp1611[57], tmp1611[56], tmp1611[55], tmp1611[54], tmp1611[53], tmp1611[52], tmp1611[51], tmp1611[50], tmp1611[49], tmp1611[48], tmp1611[47], tmp1611[46], tmp1611[45], tmp1611[44], tmp1611[43], tmp1611[42], tmp1611[41], tmp1611[40], tmp1611[39], tmp1611[38], tmp1611[37], tmp1611[36], tmp1611[35], tmp1611[34], tmp1611[33], tmp1611[32], tmp1611[31], tmp1611[30], tmp1611[29], tmp1611[28], tmp1611[27], tmp1611[26], tmp1611[25], tmp1611[24], tmp1611[23], tmp1611[22], tmp1611[21], tmp1611[20], tmp1611[19], tmp1611[18], tmp1611[17], tmp1611[16], tmp1611[15], tmp1611[14], tmp1611[13], tmp1611[12], tmp1611[11], tmp1611[10], tmp1611[9], tmp1611[8], tmp1611[7], tmp1611[6], tmp1611[5], tmp1611[4], tmp1611[3], tmp1611[2], tmp1611[1], tmp1611[0]};
    assign tmp1613 = {tmp1612[255], tmp1612[254], tmp1612[253], tmp1612[252], tmp1612[251], tmp1612[250], tmp1612[249], tmp1612[248], tmp1612[247], tmp1612[246], tmp1612[245], tmp1612[244], tmp1612[243], tmp1612[242], tmp1612[241], tmp1612[240], tmp1612[239], tmp1612[238], tmp1612[237], tmp1612[236], tmp1612[235], tmp1612[234], tmp1612[233], tmp1612[232], tmp1612[231], tmp1612[230], tmp1612[229], tmp1612[228], tmp1612[227], tmp1612[226], tmp1612[225], tmp1612[224], tmp1612[223], tmp1612[222], tmp1612[221], tmp1612[220], tmp1612[219], tmp1612[218], tmp1612[217], tmp1612[216], tmp1612[215], tmp1612[214], tmp1612[213], tmp1612[212], tmp1612[211], tmp1612[210], tmp1612[209], tmp1612[208], tmp1612[207], tmp1612[206], tmp1612[205], tmp1612[204], tmp1612[203], tmp1612[202], tmp1612[201], tmp1612[200], tmp1612[199], tmp1612[198], tmp1612[197], tmp1612[196], tmp1612[195], tmp1612[194], tmp1612[193], tmp1612[192], tmp1612[191], tmp1612[190], tmp1612[189], tmp1612[188], tmp1612[187], tmp1612[186], tmp1612[185], tmp1612[184], tmp1612[183], tmp1612[182], tmp1612[181], tmp1612[180], tmp1612[179], tmp1612[178], tmp1612[177], tmp1612[176], tmp1612[175], tmp1612[174], tmp1612[173], tmp1612[172], tmp1612[171], tmp1612[170], tmp1612[169], tmp1612[168], tmp1612[167], tmp1612[166], tmp1612[165], tmp1612[164], tmp1612[163], tmp1612[162], tmp1612[161], tmp1612[160], tmp1612[159], tmp1612[158], tmp1612[157], tmp1612[156], tmp1612[155], tmp1612[154], tmp1612[153], tmp1612[152], tmp1612[151], tmp1612[150], tmp1612[149], tmp1612[148], tmp1612[147], tmp1612[146], tmp1612[145], tmp1612[144], tmp1612[143], tmp1612[142], tmp1612[141], tmp1612[140], tmp1612[139], tmp1612[138], tmp1612[137], tmp1612[136], tmp1612[135], tmp1612[134], tmp1612[133], tmp1612[132], tmp1612[131], tmp1612[130], tmp1612[129], tmp1612[128], tmp1612[127], tmp1612[126], tmp1612[125], tmp1612[124], tmp1612[123], tmp1612[122], tmp1612[121], tmp1612[120], tmp1612[119], tmp1612[118], tmp1612[117], tmp1612[116], tmp1612[115], tmp1612[114], tmp1612[113], tmp1612[112], tmp1612[111], tmp1612[110], tmp1612[109], tmp1612[108], tmp1612[107], tmp1612[106], tmp1612[105], tmp1612[104], tmp1612[103], tmp1612[102], tmp1612[101], tmp1612[100], tmp1612[99], tmp1612[98], tmp1612[97], tmp1612[96], tmp1612[95], tmp1612[94], tmp1612[93], tmp1612[92], tmp1612[91], tmp1612[90], tmp1612[89], tmp1612[88], tmp1612[87], tmp1612[86], tmp1612[85], tmp1612[84], tmp1612[83], tmp1612[82], tmp1612[81], tmp1612[80], tmp1612[79], tmp1612[78], tmp1612[77], tmp1612[76], tmp1612[75], tmp1612[74], tmp1612[73], tmp1612[72], tmp1612[71], tmp1612[70], tmp1612[69], tmp1612[68], tmp1612[67], tmp1612[66], tmp1612[65], tmp1612[64], tmp1612[63], tmp1612[62], tmp1612[61], tmp1612[60], tmp1612[59], tmp1612[58], tmp1612[57], tmp1612[56], tmp1612[55], tmp1612[54], tmp1612[53], tmp1612[52], tmp1612[51], tmp1612[50], tmp1612[49], tmp1612[48], tmp1612[47], tmp1612[46], tmp1612[45], tmp1612[44], tmp1612[43], tmp1612[42], tmp1612[41], tmp1612[40], tmp1612[39], tmp1612[38], tmp1612[37], tmp1612[36], tmp1612[35], tmp1612[34], tmp1612[33], tmp1612[32], tmp1612[31], tmp1612[30], tmp1612[29], tmp1612[28], tmp1612[27], tmp1612[26], tmp1612[25], tmp1612[24], tmp1612[23], tmp1612[22], tmp1612[21], tmp1612[20], tmp1612[19], tmp1612[18], tmp1612[17], tmp1612[16], tmp1612[15], tmp1612[14], tmp1612[13], tmp1612[12], tmp1612[11], tmp1612[10], tmp1612[9], tmp1612[8], tmp1612[7], tmp1612[6], tmp1612[5], tmp1612[4], tmp1612[3], tmp1612[2], tmp1612[1], tmp1612[0]};
    assign tmp1614 = {const_172_0};
    assign tmp1615 = {tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614, tmp1614};
    assign tmp1616 = {tmp1615, const_172_0};
    assign tmp1617 = {tmp13[255]};
    assign tmp1618 = tmp1616 - tmp13;
    assign tmp1619 = {tmp1618[256]};
    assign tmp1620 = {tmp1616[255]};
    assign tmp1621 = ~tmp1620;
    assign tmp1622 = tmp1619 ^ tmp1621;
    assign tmp1623 = {tmp13[255]};
    assign tmp1624 = ~tmp1623;
    assign tmp1625 = tmp1622 ^ tmp1624;
    assign tmp1626 = {const_173_0};
    assign tmp1627 = {tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626, tmp1626};
    assign tmp1628 = {tmp1627, const_173_0};
    assign tmp1629 = {tmp14[255]};
    assign tmp1630 = tmp1628 - tmp14;
    assign tmp1631 = {tmp1630[256]};
    assign tmp1632 = {tmp1628[255]};
    assign tmp1633 = ~tmp1632;
    assign tmp1634 = tmp1631 ^ tmp1633;
    assign tmp1635 = {tmp14[255]};
    assign tmp1636 = ~tmp1635;
    assign tmp1637 = tmp1634 ^ tmp1636;
    assign tmp1638 = tmp1625 & tmp1637;
    assign tmp1639 = {tmp1613[255]};
    assign tmp1640 = {const_174_0};
    assign tmp1641 = {tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640, tmp1640};
    assign tmp1642 = {tmp1641, const_174_0};
    assign tmp1643 = tmp1613 - tmp1642;
    assign tmp1644 = {tmp1643[256]};
    assign tmp1645 = {tmp1613[255]};
    assign tmp1646 = ~tmp1645;
    assign tmp1647 = tmp1644 ^ tmp1646;
    assign tmp1648 = {tmp1642[255]};
    assign tmp1649 = ~tmp1648;
    assign tmp1650 = tmp1647 ^ tmp1649;
    assign tmp1651 = tmp1613 == tmp1642;
    assign tmp1652 = tmp1650 | tmp1651;
    assign tmp1653 = tmp1638 & tmp1652;
    assign tmp1654 = {tmp13[255]};
    assign tmp1655 = {const_175_0};
    assign tmp1656 = {tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655, tmp1655};
    assign tmp1657 = {tmp1656, const_175_0};
    assign tmp1658 = tmp13 - tmp1657;
    assign tmp1659 = {tmp1658[256]};
    assign tmp1660 = {tmp13[255]};
    assign tmp1661 = ~tmp1660;
    assign tmp1662 = tmp1659 ^ tmp1661;
    assign tmp1663 = {tmp1657[255]};
    assign tmp1664 = ~tmp1663;
    assign tmp1665 = tmp1662 ^ tmp1664;
    assign tmp1666 = {tmp14[255]};
    assign tmp1667 = {const_176_0};
    assign tmp1668 = {tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667, tmp1667};
    assign tmp1669 = {tmp1668, const_176_0};
    assign tmp1670 = tmp14 - tmp1669;
    assign tmp1671 = {tmp1670[256]};
    assign tmp1672 = {tmp14[255]};
    assign tmp1673 = ~tmp1672;
    assign tmp1674 = tmp1671 ^ tmp1673;
    assign tmp1675 = {tmp1669[255]};
    assign tmp1676 = ~tmp1675;
    assign tmp1677 = tmp1674 ^ tmp1676;
    assign tmp1678 = tmp1665 & tmp1677;
    assign tmp1679 = {const_177_0};
    assign tmp1680 = {tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679, tmp1679};
    assign tmp1681 = {tmp1680, const_177_0};
    assign tmp1682 = {tmp1613[255]};
    assign tmp1683 = tmp1681 - tmp1613;
    assign tmp1684 = {tmp1683[256]};
    assign tmp1685 = {tmp1681[255]};
    assign tmp1686 = ~tmp1685;
    assign tmp1687 = tmp1684 ^ tmp1686;
    assign tmp1688 = {tmp1613[255]};
    assign tmp1689 = ~tmp1688;
    assign tmp1690 = tmp1687 ^ tmp1689;
    assign tmp1691 = tmp1681 == tmp1613;
    assign tmp1692 = tmp1690 | tmp1691;
    assign tmp1693 = tmp1678 & tmp1692;
    assign tmp1694 = tmp1653 ? const_178_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp1613;
    assign tmp1695 = tmp1693 ? _ver_out_tmp_69 : tmp1694;
    assign tmp1696 = ~tmp35;
    assign tmp1697 = ~tmp36;
    assign tmp1698 = tmp1696 & tmp1697;
    assign tmp1699 = ~tmp57;
    assign tmp1700 = tmp1698 & tmp1699;
    assign tmp1701 = tmp1700 & tmp1034;
    assign tmp1702 = ~tmp1049;
    assign tmp1703 = tmp1701 & tmp1702;
    assign tmp1704 = ~tmp1050;
    assign tmp1705 = tmp1703 & tmp1704;
    assign tmp1706 = ~tmp1097;
    assign tmp1707 = tmp1705 & tmp1706;
    assign tmp1708 = ~tmp1372;
    assign tmp1709 = tmp1707 & tmp1708;
    assign tmp1710 = tmp1709 & tmp1483;
    assign tmp1711 = ~tmp35;
    assign tmp1712 = ~tmp36;
    assign tmp1713 = tmp1711 & tmp1712;
    assign tmp1714 = ~tmp57;
    assign tmp1715 = tmp1713 & tmp1714;
    assign tmp1716 = tmp1715 & tmp1034;
    assign tmp1717 = ~tmp1049;
    assign tmp1718 = tmp1716 & tmp1717;
    assign tmp1719 = ~tmp1050;
    assign tmp1720 = tmp1718 & tmp1719;
    assign tmp1721 = ~tmp1097;
    assign tmp1722 = tmp1720 & tmp1721;
    assign tmp1723 = ~tmp1372;
    assign tmp1724 = tmp1722 & tmp1723;
    assign tmp1725 = tmp1724 & tmp1483;
    assign tmp1726 = {tmp15[255]};
    assign tmp1727 = {tmp1726};
    assign tmp1728 = {tmp1727, tmp15};
    assign tmp1729 = {tmp16[255]};
    assign tmp1730 = {tmp1729};
    assign tmp1731 = {tmp1730, tmp16};
    assign tmp1732 = tmp1728 + tmp1731;
    assign tmp1733 = {tmp1732[256], tmp1732[255], tmp1732[254], tmp1732[253], tmp1732[252], tmp1732[251], tmp1732[250], tmp1732[249], tmp1732[248], tmp1732[247], tmp1732[246], tmp1732[245], tmp1732[244], tmp1732[243], tmp1732[242], tmp1732[241], tmp1732[240], tmp1732[239], tmp1732[238], tmp1732[237], tmp1732[236], tmp1732[235], tmp1732[234], tmp1732[233], tmp1732[232], tmp1732[231], tmp1732[230], tmp1732[229], tmp1732[228], tmp1732[227], tmp1732[226], tmp1732[225], tmp1732[224], tmp1732[223], tmp1732[222], tmp1732[221], tmp1732[220], tmp1732[219], tmp1732[218], tmp1732[217], tmp1732[216], tmp1732[215], tmp1732[214], tmp1732[213], tmp1732[212], tmp1732[211], tmp1732[210], tmp1732[209], tmp1732[208], tmp1732[207], tmp1732[206], tmp1732[205], tmp1732[204], tmp1732[203], tmp1732[202], tmp1732[201], tmp1732[200], tmp1732[199], tmp1732[198], tmp1732[197], tmp1732[196], tmp1732[195], tmp1732[194], tmp1732[193], tmp1732[192], tmp1732[191], tmp1732[190], tmp1732[189], tmp1732[188], tmp1732[187], tmp1732[186], tmp1732[185], tmp1732[184], tmp1732[183], tmp1732[182], tmp1732[181], tmp1732[180], tmp1732[179], tmp1732[178], tmp1732[177], tmp1732[176], tmp1732[175], tmp1732[174], tmp1732[173], tmp1732[172], tmp1732[171], tmp1732[170], tmp1732[169], tmp1732[168], tmp1732[167], tmp1732[166], tmp1732[165], tmp1732[164], tmp1732[163], tmp1732[162], tmp1732[161], tmp1732[160], tmp1732[159], tmp1732[158], tmp1732[157], tmp1732[156], tmp1732[155], tmp1732[154], tmp1732[153], tmp1732[152], tmp1732[151], tmp1732[150], tmp1732[149], tmp1732[148], tmp1732[147], tmp1732[146], tmp1732[145], tmp1732[144], tmp1732[143], tmp1732[142], tmp1732[141], tmp1732[140], tmp1732[139], tmp1732[138], tmp1732[137], tmp1732[136], tmp1732[135], tmp1732[134], tmp1732[133], tmp1732[132], tmp1732[131], tmp1732[130], tmp1732[129], tmp1732[128], tmp1732[127], tmp1732[126], tmp1732[125], tmp1732[124], tmp1732[123], tmp1732[122], tmp1732[121], tmp1732[120], tmp1732[119], tmp1732[118], tmp1732[117], tmp1732[116], tmp1732[115], tmp1732[114], tmp1732[113], tmp1732[112], tmp1732[111], tmp1732[110], tmp1732[109], tmp1732[108], tmp1732[107], tmp1732[106], tmp1732[105], tmp1732[104], tmp1732[103], tmp1732[102], tmp1732[101], tmp1732[100], tmp1732[99], tmp1732[98], tmp1732[97], tmp1732[96], tmp1732[95], tmp1732[94], tmp1732[93], tmp1732[92], tmp1732[91], tmp1732[90], tmp1732[89], tmp1732[88], tmp1732[87], tmp1732[86], tmp1732[85], tmp1732[84], tmp1732[83], tmp1732[82], tmp1732[81], tmp1732[80], tmp1732[79], tmp1732[78], tmp1732[77], tmp1732[76], tmp1732[75], tmp1732[74], tmp1732[73], tmp1732[72], tmp1732[71], tmp1732[70], tmp1732[69], tmp1732[68], tmp1732[67], tmp1732[66], tmp1732[65], tmp1732[64], tmp1732[63], tmp1732[62], tmp1732[61], tmp1732[60], tmp1732[59], tmp1732[58], tmp1732[57], tmp1732[56], tmp1732[55], tmp1732[54], tmp1732[53], tmp1732[52], tmp1732[51], tmp1732[50], tmp1732[49], tmp1732[48], tmp1732[47], tmp1732[46], tmp1732[45], tmp1732[44], tmp1732[43], tmp1732[42], tmp1732[41], tmp1732[40], tmp1732[39], tmp1732[38], tmp1732[37], tmp1732[36], tmp1732[35], tmp1732[34], tmp1732[33], tmp1732[32], tmp1732[31], tmp1732[30], tmp1732[29], tmp1732[28], tmp1732[27], tmp1732[26], tmp1732[25], tmp1732[24], tmp1732[23], tmp1732[22], tmp1732[21], tmp1732[20], tmp1732[19], tmp1732[18], tmp1732[17], tmp1732[16], tmp1732[15], tmp1732[14], tmp1732[13], tmp1732[12], tmp1732[11], tmp1732[10], tmp1732[9], tmp1732[8], tmp1732[7], tmp1732[6], tmp1732[5], tmp1732[4], tmp1732[3], tmp1732[2], tmp1732[1], tmp1732[0]};
    assign tmp1734 = {tmp1733[255], tmp1733[254], tmp1733[253], tmp1733[252], tmp1733[251], tmp1733[250], tmp1733[249], tmp1733[248], tmp1733[247], tmp1733[246], tmp1733[245], tmp1733[244], tmp1733[243], tmp1733[242], tmp1733[241], tmp1733[240], tmp1733[239], tmp1733[238], tmp1733[237], tmp1733[236], tmp1733[235], tmp1733[234], tmp1733[233], tmp1733[232], tmp1733[231], tmp1733[230], tmp1733[229], tmp1733[228], tmp1733[227], tmp1733[226], tmp1733[225], tmp1733[224], tmp1733[223], tmp1733[222], tmp1733[221], tmp1733[220], tmp1733[219], tmp1733[218], tmp1733[217], tmp1733[216], tmp1733[215], tmp1733[214], tmp1733[213], tmp1733[212], tmp1733[211], tmp1733[210], tmp1733[209], tmp1733[208], tmp1733[207], tmp1733[206], tmp1733[205], tmp1733[204], tmp1733[203], tmp1733[202], tmp1733[201], tmp1733[200], tmp1733[199], tmp1733[198], tmp1733[197], tmp1733[196], tmp1733[195], tmp1733[194], tmp1733[193], tmp1733[192], tmp1733[191], tmp1733[190], tmp1733[189], tmp1733[188], tmp1733[187], tmp1733[186], tmp1733[185], tmp1733[184], tmp1733[183], tmp1733[182], tmp1733[181], tmp1733[180], tmp1733[179], tmp1733[178], tmp1733[177], tmp1733[176], tmp1733[175], tmp1733[174], tmp1733[173], tmp1733[172], tmp1733[171], tmp1733[170], tmp1733[169], tmp1733[168], tmp1733[167], tmp1733[166], tmp1733[165], tmp1733[164], tmp1733[163], tmp1733[162], tmp1733[161], tmp1733[160], tmp1733[159], tmp1733[158], tmp1733[157], tmp1733[156], tmp1733[155], tmp1733[154], tmp1733[153], tmp1733[152], tmp1733[151], tmp1733[150], tmp1733[149], tmp1733[148], tmp1733[147], tmp1733[146], tmp1733[145], tmp1733[144], tmp1733[143], tmp1733[142], tmp1733[141], tmp1733[140], tmp1733[139], tmp1733[138], tmp1733[137], tmp1733[136], tmp1733[135], tmp1733[134], tmp1733[133], tmp1733[132], tmp1733[131], tmp1733[130], tmp1733[129], tmp1733[128], tmp1733[127], tmp1733[126], tmp1733[125], tmp1733[124], tmp1733[123], tmp1733[122], tmp1733[121], tmp1733[120], tmp1733[119], tmp1733[118], tmp1733[117], tmp1733[116], tmp1733[115], tmp1733[114], tmp1733[113], tmp1733[112], tmp1733[111], tmp1733[110], tmp1733[109], tmp1733[108], tmp1733[107], tmp1733[106], tmp1733[105], tmp1733[104], tmp1733[103], tmp1733[102], tmp1733[101], tmp1733[100], tmp1733[99], tmp1733[98], tmp1733[97], tmp1733[96], tmp1733[95], tmp1733[94], tmp1733[93], tmp1733[92], tmp1733[91], tmp1733[90], tmp1733[89], tmp1733[88], tmp1733[87], tmp1733[86], tmp1733[85], tmp1733[84], tmp1733[83], tmp1733[82], tmp1733[81], tmp1733[80], tmp1733[79], tmp1733[78], tmp1733[77], tmp1733[76], tmp1733[75], tmp1733[74], tmp1733[73], tmp1733[72], tmp1733[71], tmp1733[70], tmp1733[69], tmp1733[68], tmp1733[67], tmp1733[66], tmp1733[65], tmp1733[64], tmp1733[63], tmp1733[62], tmp1733[61], tmp1733[60], tmp1733[59], tmp1733[58], tmp1733[57], tmp1733[56], tmp1733[55], tmp1733[54], tmp1733[53], tmp1733[52], tmp1733[51], tmp1733[50], tmp1733[49], tmp1733[48], tmp1733[47], tmp1733[46], tmp1733[45], tmp1733[44], tmp1733[43], tmp1733[42], tmp1733[41], tmp1733[40], tmp1733[39], tmp1733[38], tmp1733[37], tmp1733[36], tmp1733[35], tmp1733[34], tmp1733[33], tmp1733[32], tmp1733[31], tmp1733[30], tmp1733[29], tmp1733[28], tmp1733[27], tmp1733[26], tmp1733[25], tmp1733[24], tmp1733[23], tmp1733[22], tmp1733[21], tmp1733[20], tmp1733[19], tmp1733[18], tmp1733[17], tmp1733[16], tmp1733[15], tmp1733[14], tmp1733[13], tmp1733[12], tmp1733[11], tmp1733[10], tmp1733[9], tmp1733[8], tmp1733[7], tmp1733[6], tmp1733[5], tmp1733[4], tmp1733[3], tmp1733[2], tmp1733[1], tmp1733[0]};
    assign tmp1735 = {const_180_0};
    assign tmp1736 = {tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735, tmp1735};
    assign tmp1737 = {tmp1736, const_180_0};
    assign tmp1738 = {tmp15[255]};
    assign tmp1739 = tmp1737 - tmp15;
    assign tmp1740 = {tmp1739[256]};
    assign tmp1741 = {tmp1737[255]};
    assign tmp1742 = ~tmp1741;
    assign tmp1743 = tmp1740 ^ tmp1742;
    assign tmp1744 = {tmp15[255]};
    assign tmp1745 = ~tmp1744;
    assign tmp1746 = tmp1743 ^ tmp1745;
    assign tmp1747 = {const_181_0};
    assign tmp1748 = {tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747, tmp1747};
    assign tmp1749 = {tmp1748, const_181_0};
    assign tmp1750 = {tmp16[255]};
    assign tmp1751 = tmp1749 - tmp16;
    assign tmp1752 = {tmp1751[256]};
    assign tmp1753 = {tmp1749[255]};
    assign tmp1754 = ~tmp1753;
    assign tmp1755 = tmp1752 ^ tmp1754;
    assign tmp1756 = {tmp16[255]};
    assign tmp1757 = ~tmp1756;
    assign tmp1758 = tmp1755 ^ tmp1757;
    assign tmp1759 = tmp1746 & tmp1758;
    assign tmp1760 = {tmp1734[255]};
    assign tmp1761 = {const_182_0};
    assign tmp1762 = {tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761, tmp1761};
    assign tmp1763 = {tmp1762, const_182_0};
    assign tmp1764 = tmp1734 - tmp1763;
    assign tmp1765 = {tmp1764[256]};
    assign tmp1766 = {tmp1734[255]};
    assign tmp1767 = ~tmp1766;
    assign tmp1768 = tmp1765 ^ tmp1767;
    assign tmp1769 = {tmp1763[255]};
    assign tmp1770 = ~tmp1769;
    assign tmp1771 = tmp1768 ^ tmp1770;
    assign tmp1772 = tmp1734 == tmp1763;
    assign tmp1773 = tmp1771 | tmp1772;
    assign tmp1774 = tmp1759 & tmp1773;
    assign tmp1775 = {tmp15[255]};
    assign tmp1776 = {const_183_0};
    assign tmp1777 = {tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776, tmp1776};
    assign tmp1778 = {tmp1777, const_183_0};
    assign tmp1779 = tmp15 - tmp1778;
    assign tmp1780 = {tmp1779[256]};
    assign tmp1781 = {tmp15[255]};
    assign tmp1782 = ~tmp1781;
    assign tmp1783 = tmp1780 ^ tmp1782;
    assign tmp1784 = {tmp1778[255]};
    assign tmp1785 = ~tmp1784;
    assign tmp1786 = tmp1783 ^ tmp1785;
    assign tmp1787 = {tmp16[255]};
    assign tmp1788 = {const_184_0};
    assign tmp1789 = {tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788, tmp1788};
    assign tmp1790 = {tmp1789, const_184_0};
    assign tmp1791 = tmp16 - tmp1790;
    assign tmp1792 = {tmp1791[256]};
    assign tmp1793 = {tmp16[255]};
    assign tmp1794 = ~tmp1793;
    assign tmp1795 = tmp1792 ^ tmp1794;
    assign tmp1796 = {tmp1790[255]};
    assign tmp1797 = ~tmp1796;
    assign tmp1798 = tmp1795 ^ tmp1797;
    assign tmp1799 = tmp1786 & tmp1798;
    assign tmp1800 = {const_185_0};
    assign tmp1801 = {tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800, tmp1800};
    assign tmp1802 = {tmp1801, const_185_0};
    assign tmp1803 = {tmp1734[255]};
    assign tmp1804 = tmp1802 - tmp1734;
    assign tmp1805 = {tmp1804[256]};
    assign tmp1806 = {tmp1802[255]};
    assign tmp1807 = ~tmp1806;
    assign tmp1808 = tmp1805 ^ tmp1807;
    assign tmp1809 = {tmp1734[255]};
    assign tmp1810 = ~tmp1809;
    assign tmp1811 = tmp1808 ^ tmp1810;
    assign tmp1812 = tmp1802 == tmp1734;
    assign tmp1813 = tmp1811 | tmp1812;
    assign tmp1814 = tmp1799 & tmp1813;
    assign tmp1815 = tmp1774 ? const_186_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp1734;
    assign tmp1816 = tmp1814 ? _ver_out_tmp_70 : tmp1815;
    assign tmp1817 = ~tmp35;
    assign tmp1818 = ~tmp36;
    assign tmp1819 = tmp1817 & tmp1818;
    assign tmp1820 = ~tmp57;
    assign tmp1821 = tmp1819 & tmp1820;
    assign tmp1822 = tmp1821 & tmp1034;
    assign tmp1823 = ~tmp1049;
    assign tmp1824 = tmp1822 & tmp1823;
    assign tmp1825 = ~tmp1050;
    assign tmp1826 = tmp1824 & tmp1825;
    assign tmp1827 = ~tmp1097;
    assign tmp1828 = tmp1826 & tmp1827;
    assign tmp1829 = ~tmp1372;
    assign tmp1830 = tmp1828 & tmp1829;
    assign tmp1831 = tmp1830 & tmp1483;
    assign tmp1832 = ~tmp35;
    assign tmp1833 = ~tmp36;
    assign tmp1834 = tmp1832 & tmp1833;
    assign tmp1835 = ~tmp57;
    assign tmp1836 = tmp1834 & tmp1835;
    assign tmp1837 = tmp1836 & tmp1034;
    assign tmp1838 = ~tmp1049;
    assign tmp1839 = tmp1837 & tmp1838;
    assign tmp1840 = ~tmp1050;
    assign tmp1841 = tmp1839 & tmp1840;
    assign tmp1842 = ~tmp1097;
    assign tmp1843 = tmp1841 & tmp1842;
    assign tmp1844 = ~tmp1372;
    assign tmp1845 = tmp1843 & tmp1844;
    assign tmp1846 = tmp1845 & tmp1483;
    assign tmp1847 = {tmp17[255]};
    assign tmp1848 = {tmp1847};
    assign tmp1849 = {tmp1848, tmp17};
    assign tmp1850 = {tmp18[255]};
    assign tmp1851 = {tmp1850};
    assign tmp1852 = {tmp1851, tmp18};
    assign tmp1853 = tmp1849 + tmp1852;
    assign tmp1854 = {tmp1853[256], tmp1853[255], tmp1853[254], tmp1853[253], tmp1853[252], tmp1853[251], tmp1853[250], tmp1853[249], tmp1853[248], tmp1853[247], tmp1853[246], tmp1853[245], tmp1853[244], tmp1853[243], tmp1853[242], tmp1853[241], tmp1853[240], tmp1853[239], tmp1853[238], tmp1853[237], tmp1853[236], tmp1853[235], tmp1853[234], tmp1853[233], tmp1853[232], tmp1853[231], tmp1853[230], tmp1853[229], tmp1853[228], tmp1853[227], tmp1853[226], tmp1853[225], tmp1853[224], tmp1853[223], tmp1853[222], tmp1853[221], tmp1853[220], tmp1853[219], tmp1853[218], tmp1853[217], tmp1853[216], tmp1853[215], tmp1853[214], tmp1853[213], tmp1853[212], tmp1853[211], tmp1853[210], tmp1853[209], tmp1853[208], tmp1853[207], tmp1853[206], tmp1853[205], tmp1853[204], tmp1853[203], tmp1853[202], tmp1853[201], tmp1853[200], tmp1853[199], tmp1853[198], tmp1853[197], tmp1853[196], tmp1853[195], tmp1853[194], tmp1853[193], tmp1853[192], tmp1853[191], tmp1853[190], tmp1853[189], tmp1853[188], tmp1853[187], tmp1853[186], tmp1853[185], tmp1853[184], tmp1853[183], tmp1853[182], tmp1853[181], tmp1853[180], tmp1853[179], tmp1853[178], tmp1853[177], tmp1853[176], tmp1853[175], tmp1853[174], tmp1853[173], tmp1853[172], tmp1853[171], tmp1853[170], tmp1853[169], tmp1853[168], tmp1853[167], tmp1853[166], tmp1853[165], tmp1853[164], tmp1853[163], tmp1853[162], tmp1853[161], tmp1853[160], tmp1853[159], tmp1853[158], tmp1853[157], tmp1853[156], tmp1853[155], tmp1853[154], tmp1853[153], tmp1853[152], tmp1853[151], tmp1853[150], tmp1853[149], tmp1853[148], tmp1853[147], tmp1853[146], tmp1853[145], tmp1853[144], tmp1853[143], tmp1853[142], tmp1853[141], tmp1853[140], tmp1853[139], tmp1853[138], tmp1853[137], tmp1853[136], tmp1853[135], tmp1853[134], tmp1853[133], tmp1853[132], tmp1853[131], tmp1853[130], tmp1853[129], tmp1853[128], tmp1853[127], tmp1853[126], tmp1853[125], tmp1853[124], tmp1853[123], tmp1853[122], tmp1853[121], tmp1853[120], tmp1853[119], tmp1853[118], tmp1853[117], tmp1853[116], tmp1853[115], tmp1853[114], tmp1853[113], tmp1853[112], tmp1853[111], tmp1853[110], tmp1853[109], tmp1853[108], tmp1853[107], tmp1853[106], tmp1853[105], tmp1853[104], tmp1853[103], tmp1853[102], tmp1853[101], tmp1853[100], tmp1853[99], tmp1853[98], tmp1853[97], tmp1853[96], tmp1853[95], tmp1853[94], tmp1853[93], tmp1853[92], tmp1853[91], tmp1853[90], tmp1853[89], tmp1853[88], tmp1853[87], tmp1853[86], tmp1853[85], tmp1853[84], tmp1853[83], tmp1853[82], tmp1853[81], tmp1853[80], tmp1853[79], tmp1853[78], tmp1853[77], tmp1853[76], tmp1853[75], tmp1853[74], tmp1853[73], tmp1853[72], tmp1853[71], tmp1853[70], tmp1853[69], tmp1853[68], tmp1853[67], tmp1853[66], tmp1853[65], tmp1853[64], tmp1853[63], tmp1853[62], tmp1853[61], tmp1853[60], tmp1853[59], tmp1853[58], tmp1853[57], tmp1853[56], tmp1853[55], tmp1853[54], tmp1853[53], tmp1853[52], tmp1853[51], tmp1853[50], tmp1853[49], tmp1853[48], tmp1853[47], tmp1853[46], tmp1853[45], tmp1853[44], tmp1853[43], tmp1853[42], tmp1853[41], tmp1853[40], tmp1853[39], tmp1853[38], tmp1853[37], tmp1853[36], tmp1853[35], tmp1853[34], tmp1853[33], tmp1853[32], tmp1853[31], tmp1853[30], tmp1853[29], tmp1853[28], tmp1853[27], tmp1853[26], tmp1853[25], tmp1853[24], tmp1853[23], tmp1853[22], tmp1853[21], tmp1853[20], tmp1853[19], tmp1853[18], tmp1853[17], tmp1853[16], tmp1853[15], tmp1853[14], tmp1853[13], tmp1853[12], tmp1853[11], tmp1853[10], tmp1853[9], tmp1853[8], tmp1853[7], tmp1853[6], tmp1853[5], tmp1853[4], tmp1853[3], tmp1853[2], tmp1853[1], tmp1853[0]};
    assign tmp1855 = {tmp1854[255], tmp1854[254], tmp1854[253], tmp1854[252], tmp1854[251], tmp1854[250], tmp1854[249], tmp1854[248], tmp1854[247], tmp1854[246], tmp1854[245], tmp1854[244], tmp1854[243], tmp1854[242], tmp1854[241], tmp1854[240], tmp1854[239], tmp1854[238], tmp1854[237], tmp1854[236], tmp1854[235], tmp1854[234], tmp1854[233], tmp1854[232], tmp1854[231], tmp1854[230], tmp1854[229], tmp1854[228], tmp1854[227], tmp1854[226], tmp1854[225], tmp1854[224], tmp1854[223], tmp1854[222], tmp1854[221], tmp1854[220], tmp1854[219], tmp1854[218], tmp1854[217], tmp1854[216], tmp1854[215], tmp1854[214], tmp1854[213], tmp1854[212], tmp1854[211], tmp1854[210], tmp1854[209], tmp1854[208], tmp1854[207], tmp1854[206], tmp1854[205], tmp1854[204], tmp1854[203], tmp1854[202], tmp1854[201], tmp1854[200], tmp1854[199], tmp1854[198], tmp1854[197], tmp1854[196], tmp1854[195], tmp1854[194], tmp1854[193], tmp1854[192], tmp1854[191], tmp1854[190], tmp1854[189], tmp1854[188], tmp1854[187], tmp1854[186], tmp1854[185], tmp1854[184], tmp1854[183], tmp1854[182], tmp1854[181], tmp1854[180], tmp1854[179], tmp1854[178], tmp1854[177], tmp1854[176], tmp1854[175], tmp1854[174], tmp1854[173], tmp1854[172], tmp1854[171], tmp1854[170], tmp1854[169], tmp1854[168], tmp1854[167], tmp1854[166], tmp1854[165], tmp1854[164], tmp1854[163], tmp1854[162], tmp1854[161], tmp1854[160], tmp1854[159], tmp1854[158], tmp1854[157], tmp1854[156], tmp1854[155], tmp1854[154], tmp1854[153], tmp1854[152], tmp1854[151], tmp1854[150], tmp1854[149], tmp1854[148], tmp1854[147], tmp1854[146], tmp1854[145], tmp1854[144], tmp1854[143], tmp1854[142], tmp1854[141], tmp1854[140], tmp1854[139], tmp1854[138], tmp1854[137], tmp1854[136], tmp1854[135], tmp1854[134], tmp1854[133], tmp1854[132], tmp1854[131], tmp1854[130], tmp1854[129], tmp1854[128], tmp1854[127], tmp1854[126], tmp1854[125], tmp1854[124], tmp1854[123], tmp1854[122], tmp1854[121], tmp1854[120], tmp1854[119], tmp1854[118], tmp1854[117], tmp1854[116], tmp1854[115], tmp1854[114], tmp1854[113], tmp1854[112], tmp1854[111], tmp1854[110], tmp1854[109], tmp1854[108], tmp1854[107], tmp1854[106], tmp1854[105], tmp1854[104], tmp1854[103], tmp1854[102], tmp1854[101], tmp1854[100], tmp1854[99], tmp1854[98], tmp1854[97], tmp1854[96], tmp1854[95], tmp1854[94], tmp1854[93], tmp1854[92], tmp1854[91], tmp1854[90], tmp1854[89], tmp1854[88], tmp1854[87], tmp1854[86], tmp1854[85], tmp1854[84], tmp1854[83], tmp1854[82], tmp1854[81], tmp1854[80], tmp1854[79], tmp1854[78], tmp1854[77], tmp1854[76], tmp1854[75], tmp1854[74], tmp1854[73], tmp1854[72], tmp1854[71], tmp1854[70], tmp1854[69], tmp1854[68], tmp1854[67], tmp1854[66], tmp1854[65], tmp1854[64], tmp1854[63], tmp1854[62], tmp1854[61], tmp1854[60], tmp1854[59], tmp1854[58], tmp1854[57], tmp1854[56], tmp1854[55], tmp1854[54], tmp1854[53], tmp1854[52], tmp1854[51], tmp1854[50], tmp1854[49], tmp1854[48], tmp1854[47], tmp1854[46], tmp1854[45], tmp1854[44], tmp1854[43], tmp1854[42], tmp1854[41], tmp1854[40], tmp1854[39], tmp1854[38], tmp1854[37], tmp1854[36], tmp1854[35], tmp1854[34], tmp1854[33], tmp1854[32], tmp1854[31], tmp1854[30], tmp1854[29], tmp1854[28], tmp1854[27], tmp1854[26], tmp1854[25], tmp1854[24], tmp1854[23], tmp1854[22], tmp1854[21], tmp1854[20], tmp1854[19], tmp1854[18], tmp1854[17], tmp1854[16], tmp1854[15], tmp1854[14], tmp1854[13], tmp1854[12], tmp1854[11], tmp1854[10], tmp1854[9], tmp1854[8], tmp1854[7], tmp1854[6], tmp1854[5], tmp1854[4], tmp1854[3], tmp1854[2], tmp1854[1], tmp1854[0]};
    assign tmp1856 = {const_188_0};
    assign tmp1857 = {tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856, tmp1856};
    assign tmp1858 = {tmp1857, const_188_0};
    assign tmp1859 = {tmp17[255]};
    assign tmp1860 = tmp1858 - tmp17;
    assign tmp1861 = {tmp1860[256]};
    assign tmp1862 = {tmp1858[255]};
    assign tmp1863 = ~tmp1862;
    assign tmp1864 = tmp1861 ^ tmp1863;
    assign tmp1865 = {tmp17[255]};
    assign tmp1866 = ~tmp1865;
    assign tmp1867 = tmp1864 ^ tmp1866;
    assign tmp1868 = {const_189_0};
    assign tmp1869 = {tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868, tmp1868};
    assign tmp1870 = {tmp1869, const_189_0};
    assign tmp1871 = {tmp18[255]};
    assign tmp1872 = tmp1870 - tmp18;
    assign tmp1873 = {tmp1872[256]};
    assign tmp1874 = {tmp1870[255]};
    assign tmp1875 = ~tmp1874;
    assign tmp1876 = tmp1873 ^ tmp1875;
    assign tmp1877 = {tmp18[255]};
    assign tmp1878 = ~tmp1877;
    assign tmp1879 = tmp1876 ^ tmp1878;
    assign tmp1880 = tmp1867 & tmp1879;
    assign tmp1881 = {tmp1855[255]};
    assign tmp1882 = {const_190_0};
    assign tmp1883 = {tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882, tmp1882};
    assign tmp1884 = {tmp1883, const_190_0};
    assign tmp1885 = tmp1855 - tmp1884;
    assign tmp1886 = {tmp1885[256]};
    assign tmp1887 = {tmp1855[255]};
    assign tmp1888 = ~tmp1887;
    assign tmp1889 = tmp1886 ^ tmp1888;
    assign tmp1890 = {tmp1884[255]};
    assign tmp1891 = ~tmp1890;
    assign tmp1892 = tmp1889 ^ tmp1891;
    assign tmp1893 = tmp1855 == tmp1884;
    assign tmp1894 = tmp1892 | tmp1893;
    assign tmp1895 = tmp1880 & tmp1894;
    assign tmp1896 = {tmp17[255]};
    assign tmp1897 = {const_191_0};
    assign tmp1898 = {tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897, tmp1897};
    assign tmp1899 = {tmp1898, const_191_0};
    assign tmp1900 = tmp17 - tmp1899;
    assign tmp1901 = {tmp1900[256]};
    assign tmp1902 = {tmp17[255]};
    assign tmp1903 = ~tmp1902;
    assign tmp1904 = tmp1901 ^ tmp1903;
    assign tmp1905 = {tmp1899[255]};
    assign tmp1906 = ~tmp1905;
    assign tmp1907 = tmp1904 ^ tmp1906;
    assign tmp1908 = {tmp18[255]};
    assign tmp1909 = {const_192_0};
    assign tmp1910 = {tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909, tmp1909};
    assign tmp1911 = {tmp1910, const_192_0};
    assign tmp1912 = tmp18 - tmp1911;
    assign tmp1913 = {tmp1912[256]};
    assign tmp1914 = {tmp18[255]};
    assign tmp1915 = ~tmp1914;
    assign tmp1916 = tmp1913 ^ tmp1915;
    assign tmp1917 = {tmp1911[255]};
    assign tmp1918 = ~tmp1917;
    assign tmp1919 = tmp1916 ^ tmp1918;
    assign tmp1920 = tmp1907 & tmp1919;
    assign tmp1921 = {const_193_0};
    assign tmp1922 = {tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921, tmp1921};
    assign tmp1923 = {tmp1922, const_193_0};
    assign tmp1924 = {tmp1855[255]};
    assign tmp1925 = tmp1923 - tmp1855;
    assign tmp1926 = {tmp1925[256]};
    assign tmp1927 = {tmp1923[255]};
    assign tmp1928 = ~tmp1927;
    assign tmp1929 = tmp1926 ^ tmp1928;
    assign tmp1930 = {tmp1855[255]};
    assign tmp1931 = ~tmp1930;
    assign tmp1932 = tmp1929 ^ tmp1931;
    assign tmp1933 = tmp1923 == tmp1855;
    assign tmp1934 = tmp1932 | tmp1933;
    assign tmp1935 = tmp1920 & tmp1934;
    assign tmp1936 = tmp1895 ? const_194_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp1855;
    assign tmp1937 = tmp1935 ? _ver_out_tmp_73 : tmp1936;
    assign tmp1938 = ~tmp35;
    assign tmp1939 = ~tmp36;
    assign tmp1940 = tmp1938 & tmp1939;
    assign tmp1941 = ~tmp57;
    assign tmp1942 = tmp1940 & tmp1941;
    assign tmp1943 = tmp1942 & tmp1034;
    assign tmp1944 = ~tmp1049;
    assign tmp1945 = tmp1943 & tmp1944;
    assign tmp1946 = ~tmp1050;
    assign tmp1947 = tmp1945 & tmp1946;
    assign tmp1948 = ~tmp1097;
    assign tmp1949 = tmp1947 & tmp1948;
    assign tmp1950 = ~tmp1372;
    assign tmp1951 = tmp1949 & tmp1950;
    assign tmp1952 = tmp1951 & tmp1483;
    assign tmp1953 = ~tmp35;
    assign tmp1954 = ~tmp36;
    assign tmp1955 = tmp1953 & tmp1954;
    assign tmp1956 = ~tmp57;
    assign tmp1957 = tmp1955 & tmp1956;
    assign tmp1958 = tmp1957 & tmp1034;
    assign tmp1959 = ~tmp1049;
    assign tmp1960 = tmp1958 & tmp1959;
    assign tmp1961 = ~tmp1050;
    assign tmp1962 = tmp1960 & tmp1961;
    assign tmp1963 = ~tmp1097;
    assign tmp1964 = tmp1962 & tmp1963;
    assign tmp1965 = ~tmp1372;
    assign tmp1966 = tmp1964 & tmp1965;
    assign tmp1967 = tmp1966 & tmp1483;
    assign tmp1968 = my_calculator_in_y == const_196_8;
    assign tmp1969 = tmp11 == _ver_out_tmp_74;
    assign tmp1970 = {const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0, const_199_0};
    assign tmp1971 = {tmp1970, const_198_0};
    assign tmp1972 = tmp1971 - tmp11;
    assign tmp1973 = {const_201_0, const_201_0};
    assign tmp1974 = {tmp1973, const_200_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp1975 = tmp1969 ? tmp1974 : tmp1972;
    assign tmp1976 = {tmp1975[255], tmp1975[254], tmp1975[253], tmp1975[252], tmp1975[251], tmp1975[250], tmp1975[249], tmp1975[248], tmp1975[247], tmp1975[246], tmp1975[245], tmp1975[244], tmp1975[243], tmp1975[242], tmp1975[241], tmp1975[240], tmp1975[239], tmp1975[238], tmp1975[237], tmp1975[236], tmp1975[235], tmp1975[234], tmp1975[233], tmp1975[232], tmp1975[231], tmp1975[230], tmp1975[229], tmp1975[228], tmp1975[227], tmp1975[226], tmp1975[225], tmp1975[224], tmp1975[223], tmp1975[222], tmp1975[221], tmp1975[220], tmp1975[219], tmp1975[218], tmp1975[217], tmp1975[216], tmp1975[215], tmp1975[214], tmp1975[213], tmp1975[212], tmp1975[211], tmp1975[210], tmp1975[209], tmp1975[208], tmp1975[207], tmp1975[206], tmp1975[205], tmp1975[204], tmp1975[203], tmp1975[202], tmp1975[201], tmp1975[200], tmp1975[199], tmp1975[198], tmp1975[197], tmp1975[196], tmp1975[195], tmp1975[194], tmp1975[193], tmp1975[192], tmp1975[191], tmp1975[190], tmp1975[189], tmp1975[188], tmp1975[187], tmp1975[186], tmp1975[185], tmp1975[184], tmp1975[183], tmp1975[182], tmp1975[181], tmp1975[180], tmp1975[179], tmp1975[178], tmp1975[177], tmp1975[176], tmp1975[175], tmp1975[174], tmp1975[173], tmp1975[172], tmp1975[171], tmp1975[170], tmp1975[169], tmp1975[168], tmp1975[167], tmp1975[166], tmp1975[165], tmp1975[164], tmp1975[163], tmp1975[162], tmp1975[161], tmp1975[160], tmp1975[159], tmp1975[158], tmp1975[157], tmp1975[156], tmp1975[155], tmp1975[154], tmp1975[153], tmp1975[152], tmp1975[151], tmp1975[150], tmp1975[149], tmp1975[148], tmp1975[147], tmp1975[146], tmp1975[145], tmp1975[144], tmp1975[143], tmp1975[142], tmp1975[141], tmp1975[140], tmp1975[139], tmp1975[138], tmp1975[137], tmp1975[136], tmp1975[135], tmp1975[134], tmp1975[133], tmp1975[132], tmp1975[131], tmp1975[130], tmp1975[129], tmp1975[128], tmp1975[127], tmp1975[126], tmp1975[125], tmp1975[124], tmp1975[123], tmp1975[122], tmp1975[121], tmp1975[120], tmp1975[119], tmp1975[118], tmp1975[117], tmp1975[116], tmp1975[115], tmp1975[114], tmp1975[113], tmp1975[112], tmp1975[111], tmp1975[110], tmp1975[109], tmp1975[108], tmp1975[107], tmp1975[106], tmp1975[105], tmp1975[104], tmp1975[103], tmp1975[102], tmp1975[101], tmp1975[100], tmp1975[99], tmp1975[98], tmp1975[97], tmp1975[96], tmp1975[95], tmp1975[94], tmp1975[93], tmp1975[92], tmp1975[91], tmp1975[90], tmp1975[89], tmp1975[88], tmp1975[87], tmp1975[86], tmp1975[85], tmp1975[84], tmp1975[83], tmp1975[82], tmp1975[81], tmp1975[80], tmp1975[79], tmp1975[78], tmp1975[77], tmp1975[76], tmp1975[75], tmp1975[74], tmp1975[73], tmp1975[72], tmp1975[71], tmp1975[70], tmp1975[69], tmp1975[68], tmp1975[67], tmp1975[66], tmp1975[65], tmp1975[64], tmp1975[63], tmp1975[62], tmp1975[61], tmp1975[60], tmp1975[59], tmp1975[58], tmp1975[57], tmp1975[56], tmp1975[55], tmp1975[54], tmp1975[53], tmp1975[52], tmp1975[51], tmp1975[50], tmp1975[49], tmp1975[48], tmp1975[47], tmp1975[46], tmp1975[45], tmp1975[44], tmp1975[43], tmp1975[42], tmp1975[41], tmp1975[40], tmp1975[39], tmp1975[38], tmp1975[37], tmp1975[36], tmp1975[35], tmp1975[34], tmp1975[33], tmp1975[32], tmp1975[31], tmp1975[30], tmp1975[29], tmp1975[28], tmp1975[27], tmp1975[26], tmp1975[25], tmp1975[24], tmp1975[23], tmp1975[22], tmp1975[21], tmp1975[20], tmp1975[19], tmp1975[18], tmp1975[17], tmp1975[16], tmp1975[15], tmp1975[14], tmp1975[13], tmp1975[12], tmp1975[11], tmp1975[10], tmp1975[9], tmp1975[8], tmp1975[7], tmp1975[6], tmp1975[5], tmp1975[4], tmp1975[3], tmp1975[2], tmp1975[1], tmp1975[0]};
    assign tmp1977 = ~tmp35;
    assign tmp1978 = ~tmp36;
    assign tmp1979 = tmp1977 & tmp1978;
    assign tmp1980 = ~tmp57;
    assign tmp1981 = tmp1979 & tmp1980;
    assign tmp1982 = tmp1981 & tmp1034;
    assign tmp1983 = ~tmp1049;
    assign tmp1984 = tmp1982 & tmp1983;
    assign tmp1985 = ~tmp1050;
    assign tmp1986 = tmp1984 & tmp1985;
    assign tmp1987 = ~tmp1097;
    assign tmp1988 = tmp1986 & tmp1987;
    assign tmp1989 = ~tmp1372;
    assign tmp1990 = tmp1988 & tmp1989;
    assign tmp1991 = ~tmp1483;
    assign tmp1992 = tmp1990 & tmp1991;
    assign tmp1993 = tmp1992 & tmp1968;
    assign tmp1994 = tmp13 == _ver_out_tmp_76;
    assign tmp1995 = {const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0, const_204_0};
    assign tmp1996 = {tmp1995, const_203_0};
    assign tmp1997 = tmp1996 - tmp13;
    assign tmp1998 = {const_206_0, const_206_0};
    assign tmp1999 = {tmp1998, const_205_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp2000 = tmp1994 ? tmp1999 : tmp1997;
    assign tmp2001 = {tmp2000[255], tmp2000[254], tmp2000[253], tmp2000[252], tmp2000[251], tmp2000[250], tmp2000[249], tmp2000[248], tmp2000[247], tmp2000[246], tmp2000[245], tmp2000[244], tmp2000[243], tmp2000[242], tmp2000[241], tmp2000[240], tmp2000[239], tmp2000[238], tmp2000[237], tmp2000[236], tmp2000[235], tmp2000[234], tmp2000[233], tmp2000[232], tmp2000[231], tmp2000[230], tmp2000[229], tmp2000[228], tmp2000[227], tmp2000[226], tmp2000[225], tmp2000[224], tmp2000[223], tmp2000[222], tmp2000[221], tmp2000[220], tmp2000[219], tmp2000[218], tmp2000[217], tmp2000[216], tmp2000[215], tmp2000[214], tmp2000[213], tmp2000[212], tmp2000[211], tmp2000[210], tmp2000[209], tmp2000[208], tmp2000[207], tmp2000[206], tmp2000[205], tmp2000[204], tmp2000[203], tmp2000[202], tmp2000[201], tmp2000[200], tmp2000[199], tmp2000[198], tmp2000[197], tmp2000[196], tmp2000[195], tmp2000[194], tmp2000[193], tmp2000[192], tmp2000[191], tmp2000[190], tmp2000[189], tmp2000[188], tmp2000[187], tmp2000[186], tmp2000[185], tmp2000[184], tmp2000[183], tmp2000[182], tmp2000[181], tmp2000[180], tmp2000[179], tmp2000[178], tmp2000[177], tmp2000[176], tmp2000[175], tmp2000[174], tmp2000[173], tmp2000[172], tmp2000[171], tmp2000[170], tmp2000[169], tmp2000[168], tmp2000[167], tmp2000[166], tmp2000[165], tmp2000[164], tmp2000[163], tmp2000[162], tmp2000[161], tmp2000[160], tmp2000[159], tmp2000[158], tmp2000[157], tmp2000[156], tmp2000[155], tmp2000[154], tmp2000[153], tmp2000[152], tmp2000[151], tmp2000[150], tmp2000[149], tmp2000[148], tmp2000[147], tmp2000[146], tmp2000[145], tmp2000[144], tmp2000[143], tmp2000[142], tmp2000[141], tmp2000[140], tmp2000[139], tmp2000[138], tmp2000[137], tmp2000[136], tmp2000[135], tmp2000[134], tmp2000[133], tmp2000[132], tmp2000[131], tmp2000[130], tmp2000[129], tmp2000[128], tmp2000[127], tmp2000[126], tmp2000[125], tmp2000[124], tmp2000[123], tmp2000[122], tmp2000[121], tmp2000[120], tmp2000[119], tmp2000[118], tmp2000[117], tmp2000[116], tmp2000[115], tmp2000[114], tmp2000[113], tmp2000[112], tmp2000[111], tmp2000[110], tmp2000[109], tmp2000[108], tmp2000[107], tmp2000[106], tmp2000[105], tmp2000[104], tmp2000[103], tmp2000[102], tmp2000[101], tmp2000[100], tmp2000[99], tmp2000[98], tmp2000[97], tmp2000[96], tmp2000[95], tmp2000[94], tmp2000[93], tmp2000[92], tmp2000[91], tmp2000[90], tmp2000[89], tmp2000[88], tmp2000[87], tmp2000[86], tmp2000[85], tmp2000[84], tmp2000[83], tmp2000[82], tmp2000[81], tmp2000[80], tmp2000[79], tmp2000[78], tmp2000[77], tmp2000[76], tmp2000[75], tmp2000[74], tmp2000[73], tmp2000[72], tmp2000[71], tmp2000[70], tmp2000[69], tmp2000[68], tmp2000[67], tmp2000[66], tmp2000[65], tmp2000[64], tmp2000[63], tmp2000[62], tmp2000[61], tmp2000[60], tmp2000[59], tmp2000[58], tmp2000[57], tmp2000[56], tmp2000[55], tmp2000[54], tmp2000[53], tmp2000[52], tmp2000[51], tmp2000[50], tmp2000[49], tmp2000[48], tmp2000[47], tmp2000[46], tmp2000[45], tmp2000[44], tmp2000[43], tmp2000[42], tmp2000[41], tmp2000[40], tmp2000[39], tmp2000[38], tmp2000[37], tmp2000[36], tmp2000[35], tmp2000[34], tmp2000[33], tmp2000[32], tmp2000[31], tmp2000[30], tmp2000[29], tmp2000[28], tmp2000[27], tmp2000[26], tmp2000[25], tmp2000[24], tmp2000[23], tmp2000[22], tmp2000[21], tmp2000[20], tmp2000[19], tmp2000[18], tmp2000[17], tmp2000[16], tmp2000[15], tmp2000[14], tmp2000[13], tmp2000[12], tmp2000[11], tmp2000[10], tmp2000[9], tmp2000[8], tmp2000[7], tmp2000[6], tmp2000[5], tmp2000[4], tmp2000[3], tmp2000[2], tmp2000[1], tmp2000[0]};
    assign tmp2002 = ~tmp35;
    assign tmp2003 = ~tmp36;
    assign tmp2004 = tmp2002 & tmp2003;
    assign tmp2005 = ~tmp57;
    assign tmp2006 = tmp2004 & tmp2005;
    assign tmp2007 = tmp2006 & tmp1034;
    assign tmp2008 = ~tmp1049;
    assign tmp2009 = tmp2007 & tmp2008;
    assign tmp2010 = ~tmp1050;
    assign tmp2011 = tmp2009 & tmp2010;
    assign tmp2012 = ~tmp1097;
    assign tmp2013 = tmp2011 & tmp2012;
    assign tmp2014 = ~tmp1372;
    assign tmp2015 = tmp2013 & tmp2014;
    assign tmp2016 = ~tmp1483;
    assign tmp2017 = tmp2015 & tmp2016;
    assign tmp2018 = tmp2017 & tmp1968;
    assign tmp2019 = tmp15 == _ver_out_tmp_77;
    assign tmp2020 = {const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0, const_209_0};
    assign tmp2021 = {tmp2020, const_208_0};
    assign tmp2022 = tmp2021 - tmp15;
    assign tmp2023 = {const_211_0, const_211_0};
    assign tmp2024 = {tmp2023, const_210_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp2025 = tmp2019 ? tmp2024 : tmp2022;
    assign tmp2026 = {tmp2025[255], tmp2025[254], tmp2025[253], tmp2025[252], tmp2025[251], tmp2025[250], tmp2025[249], tmp2025[248], tmp2025[247], tmp2025[246], tmp2025[245], tmp2025[244], tmp2025[243], tmp2025[242], tmp2025[241], tmp2025[240], tmp2025[239], tmp2025[238], tmp2025[237], tmp2025[236], tmp2025[235], tmp2025[234], tmp2025[233], tmp2025[232], tmp2025[231], tmp2025[230], tmp2025[229], tmp2025[228], tmp2025[227], tmp2025[226], tmp2025[225], tmp2025[224], tmp2025[223], tmp2025[222], tmp2025[221], tmp2025[220], tmp2025[219], tmp2025[218], tmp2025[217], tmp2025[216], tmp2025[215], tmp2025[214], tmp2025[213], tmp2025[212], tmp2025[211], tmp2025[210], tmp2025[209], tmp2025[208], tmp2025[207], tmp2025[206], tmp2025[205], tmp2025[204], tmp2025[203], tmp2025[202], tmp2025[201], tmp2025[200], tmp2025[199], tmp2025[198], tmp2025[197], tmp2025[196], tmp2025[195], tmp2025[194], tmp2025[193], tmp2025[192], tmp2025[191], tmp2025[190], tmp2025[189], tmp2025[188], tmp2025[187], tmp2025[186], tmp2025[185], tmp2025[184], tmp2025[183], tmp2025[182], tmp2025[181], tmp2025[180], tmp2025[179], tmp2025[178], tmp2025[177], tmp2025[176], tmp2025[175], tmp2025[174], tmp2025[173], tmp2025[172], tmp2025[171], tmp2025[170], tmp2025[169], tmp2025[168], tmp2025[167], tmp2025[166], tmp2025[165], tmp2025[164], tmp2025[163], tmp2025[162], tmp2025[161], tmp2025[160], tmp2025[159], tmp2025[158], tmp2025[157], tmp2025[156], tmp2025[155], tmp2025[154], tmp2025[153], tmp2025[152], tmp2025[151], tmp2025[150], tmp2025[149], tmp2025[148], tmp2025[147], tmp2025[146], tmp2025[145], tmp2025[144], tmp2025[143], tmp2025[142], tmp2025[141], tmp2025[140], tmp2025[139], tmp2025[138], tmp2025[137], tmp2025[136], tmp2025[135], tmp2025[134], tmp2025[133], tmp2025[132], tmp2025[131], tmp2025[130], tmp2025[129], tmp2025[128], tmp2025[127], tmp2025[126], tmp2025[125], tmp2025[124], tmp2025[123], tmp2025[122], tmp2025[121], tmp2025[120], tmp2025[119], tmp2025[118], tmp2025[117], tmp2025[116], tmp2025[115], tmp2025[114], tmp2025[113], tmp2025[112], tmp2025[111], tmp2025[110], tmp2025[109], tmp2025[108], tmp2025[107], tmp2025[106], tmp2025[105], tmp2025[104], tmp2025[103], tmp2025[102], tmp2025[101], tmp2025[100], tmp2025[99], tmp2025[98], tmp2025[97], tmp2025[96], tmp2025[95], tmp2025[94], tmp2025[93], tmp2025[92], tmp2025[91], tmp2025[90], tmp2025[89], tmp2025[88], tmp2025[87], tmp2025[86], tmp2025[85], tmp2025[84], tmp2025[83], tmp2025[82], tmp2025[81], tmp2025[80], tmp2025[79], tmp2025[78], tmp2025[77], tmp2025[76], tmp2025[75], tmp2025[74], tmp2025[73], tmp2025[72], tmp2025[71], tmp2025[70], tmp2025[69], tmp2025[68], tmp2025[67], tmp2025[66], tmp2025[65], tmp2025[64], tmp2025[63], tmp2025[62], tmp2025[61], tmp2025[60], tmp2025[59], tmp2025[58], tmp2025[57], tmp2025[56], tmp2025[55], tmp2025[54], tmp2025[53], tmp2025[52], tmp2025[51], tmp2025[50], tmp2025[49], tmp2025[48], tmp2025[47], tmp2025[46], tmp2025[45], tmp2025[44], tmp2025[43], tmp2025[42], tmp2025[41], tmp2025[40], tmp2025[39], tmp2025[38], tmp2025[37], tmp2025[36], tmp2025[35], tmp2025[34], tmp2025[33], tmp2025[32], tmp2025[31], tmp2025[30], tmp2025[29], tmp2025[28], tmp2025[27], tmp2025[26], tmp2025[25], tmp2025[24], tmp2025[23], tmp2025[22], tmp2025[21], tmp2025[20], tmp2025[19], tmp2025[18], tmp2025[17], tmp2025[16], tmp2025[15], tmp2025[14], tmp2025[13], tmp2025[12], tmp2025[11], tmp2025[10], tmp2025[9], tmp2025[8], tmp2025[7], tmp2025[6], tmp2025[5], tmp2025[4], tmp2025[3], tmp2025[2], tmp2025[1], tmp2025[0]};
    assign tmp2027 = ~tmp35;
    assign tmp2028 = ~tmp36;
    assign tmp2029 = tmp2027 & tmp2028;
    assign tmp2030 = ~tmp57;
    assign tmp2031 = tmp2029 & tmp2030;
    assign tmp2032 = tmp2031 & tmp1034;
    assign tmp2033 = ~tmp1049;
    assign tmp2034 = tmp2032 & tmp2033;
    assign tmp2035 = ~tmp1050;
    assign tmp2036 = tmp2034 & tmp2035;
    assign tmp2037 = ~tmp1097;
    assign tmp2038 = tmp2036 & tmp2037;
    assign tmp2039 = ~tmp1372;
    assign tmp2040 = tmp2038 & tmp2039;
    assign tmp2041 = ~tmp1483;
    assign tmp2042 = tmp2040 & tmp2041;
    assign tmp2043 = tmp2042 & tmp1968;
    assign tmp2044 = tmp17 == _ver_out_tmp_78;
    assign tmp2045 = {const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0, const_214_0};
    assign tmp2046 = {tmp2045, const_213_0};
    assign tmp2047 = tmp2046 - tmp17;
    assign tmp2048 = {const_216_0, const_216_0};
    assign tmp2049 = {tmp2048, const_215_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp2050 = tmp2044 ? tmp2049 : tmp2047;
    assign tmp2051 = {tmp2050[255], tmp2050[254], tmp2050[253], tmp2050[252], tmp2050[251], tmp2050[250], tmp2050[249], tmp2050[248], tmp2050[247], tmp2050[246], tmp2050[245], tmp2050[244], tmp2050[243], tmp2050[242], tmp2050[241], tmp2050[240], tmp2050[239], tmp2050[238], tmp2050[237], tmp2050[236], tmp2050[235], tmp2050[234], tmp2050[233], tmp2050[232], tmp2050[231], tmp2050[230], tmp2050[229], tmp2050[228], tmp2050[227], tmp2050[226], tmp2050[225], tmp2050[224], tmp2050[223], tmp2050[222], tmp2050[221], tmp2050[220], tmp2050[219], tmp2050[218], tmp2050[217], tmp2050[216], tmp2050[215], tmp2050[214], tmp2050[213], tmp2050[212], tmp2050[211], tmp2050[210], tmp2050[209], tmp2050[208], tmp2050[207], tmp2050[206], tmp2050[205], tmp2050[204], tmp2050[203], tmp2050[202], tmp2050[201], tmp2050[200], tmp2050[199], tmp2050[198], tmp2050[197], tmp2050[196], tmp2050[195], tmp2050[194], tmp2050[193], tmp2050[192], tmp2050[191], tmp2050[190], tmp2050[189], tmp2050[188], tmp2050[187], tmp2050[186], tmp2050[185], tmp2050[184], tmp2050[183], tmp2050[182], tmp2050[181], tmp2050[180], tmp2050[179], tmp2050[178], tmp2050[177], tmp2050[176], tmp2050[175], tmp2050[174], tmp2050[173], tmp2050[172], tmp2050[171], tmp2050[170], tmp2050[169], tmp2050[168], tmp2050[167], tmp2050[166], tmp2050[165], tmp2050[164], tmp2050[163], tmp2050[162], tmp2050[161], tmp2050[160], tmp2050[159], tmp2050[158], tmp2050[157], tmp2050[156], tmp2050[155], tmp2050[154], tmp2050[153], tmp2050[152], tmp2050[151], tmp2050[150], tmp2050[149], tmp2050[148], tmp2050[147], tmp2050[146], tmp2050[145], tmp2050[144], tmp2050[143], tmp2050[142], tmp2050[141], tmp2050[140], tmp2050[139], tmp2050[138], tmp2050[137], tmp2050[136], tmp2050[135], tmp2050[134], tmp2050[133], tmp2050[132], tmp2050[131], tmp2050[130], tmp2050[129], tmp2050[128], tmp2050[127], tmp2050[126], tmp2050[125], tmp2050[124], tmp2050[123], tmp2050[122], tmp2050[121], tmp2050[120], tmp2050[119], tmp2050[118], tmp2050[117], tmp2050[116], tmp2050[115], tmp2050[114], tmp2050[113], tmp2050[112], tmp2050[111], tmp2050[110], tmp2050[109], tmp2050[108], tmp2050[107], tmp2050[106], tmp2050[105], tmp2050[104], tmp2050[103], tmp2050[102], tmp2050[101], tmp2050[100], tmp2050[99], tmp2050[98], tmp2050[97], tmp2050[96], tmp2050[95], tmp2050[94], tmp2050[93], tmp2050[92], tmp2050[91], tmp2050[90], tmp2050[89], tmp2050[88], tmp2050[87], tmp2050[86], tmp2050[85], tmp2050[84], tmp2050[83], tmp2050[82], tmp2050[81], tmp2050[80], tmp2050[79], tmp2050[78], tmp2050[77], tmp2050[76], tmp2050[75], tmp2050[74], tmp2050[73], tmp2050[72], tmp2050[71], tmp2050[70], tmp2050[69], tmp2050[68], tmp2050[67], tmp2050[66], tmp2050[65], tmp2050[64], tmp2050[63], tmp2050[62], tmp2050[61], tmp2050[60], tmp2050[59], tmp2050[58], tmp2050[57], tmp2050[56], tmp2050[55], tmp2050[54], tmp2050[53], tmp2050[52], tmp2050[51], tmp2050[50], tmp2050[49], tmp2050[48], tmp2050[47], tmp2050[46], tmp2050[45], tmp2050[44], tmp2050[43], tmp2050[42], tmp2050[41], tmp2050[40], tmp2050[39], tmp2050[38], tmp2050[37], tmp2050[36], tmp2050[35], tmp2050[34], tmp2050[33], tmp2050[32], tmp2050[31], tmp2050[30], tmp2050[29], tmp2050[28], tmp2050[27], tmp2050[26], tmp2050[25], tmp2050[24], tmp2050[23], tmp2050[22], tmp2050[21], tmp2050[20], tmp2050[19], tmp2050[18], tmp2050[17], tmp2050[16], tmp2050[15], tmp2050[14], tmp2050[13], tmp2050[12], tmp2050[11], tmp2050[10], tmp2050[9], tmp2050[8], tmp2050[7], tmp2050[6], tmp2050[5], tmp2050[4], tmp2050[3], tmp2050[2], tmp2050[1], tmp2050[0]};
    assign tmp2052 = ~tmp35;
    assign tmp2053 = ~tmp36;
    assign tmp2054 = tmp2052 & tmp2053;
    assign tmp2055 = ~tmp57;
    assign tmp2056 = tmp2054 & tmp2055;
    assign tmp2057 = tmp2056 & tmp1034;
    assign tmp2058 = ~tmp1049;
    assign tmp2059 = tmp2057 & tmp2058;
    assign tmp2060 = ~tmp1050;
    assign tmp2061 = tmp2059 & tmp2060;
    assign tmp2062 = ~tmp1097;
    assign tmp2063 = tmp2061 & tmp2062;
    assign tmp2064 = ~tmp1372;
    assign tmp2065 = tmp2063 & tmp2064;
    assign tmp2066 = ~tmp1483;
    assign tmp2067 = tmp2065 & tmp2066;
    assign tmp2068 = tmp2067 & tmp1968;
    assign tmp2069 = {const_218_0};
    assign tmp2070 = {tmp2069, const_217_3};
    assign tmp2071 = my_calculator_ctrl == tmp2070;
    assign tmp2072 = {tmp11[255]};
    assign tmp2073 = {const_219_0};
    assign tmp2074 = {tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073, tmp2073};
    assign tmp2075 = {tmp2074, const_219_0};
    assign tmp2076 = tmp11 - tmp2075;
    assign tmp2077 = {tmp2076[256]};
    assign tmp2078 = {tmp11[255]};
    assign tmp2079 = ~tmp2078;
    assign tmp2080 = tmp2077 ^ tmp2079;
    assign tmp2081 = {tmp2075[255]};
    assign tmp2082 = ~tmp2081;
    assign tmp2083 = tmp2080 ^ tmp2082;
    assign tmp2084 = {tmp12[255]};
    assign tmp2085 = {const_220_0};
    assign tmp2086 = {tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085, tmp2085};
    assign tmp2087 = {tmp2086, const_220_0};
    assign tmp2088 = tmp12 - tmp2087;
    assign tmp2089 = {tmp2088[256]};
    assign tmp2090 = {tmp12[255]};
    assign tmp2091 = ~tmp2090;
    assign tmp2092 = tmp2089 ^ tmp2091;
    assign tmp2093 = {tmp2087[255]};
    assign tmp2094 = ~tmp2093;
    assign tmp2095 = tmp2092 ^ tmp2094;
    assign tmp2096 = tmp2083 == tmp2095;
    assign tmp2097 = {tmp12[255]};
    assign tmp2098 = {const_221_0};
    assign tmp2099 = {tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098, tmp2098};
    assign tmp2100 = {tmp2099, const_221_0};
    assign tmp2101 = tmp12 - tmp2100;
    assign tmp2102 = {tmp2101[256]};
    assign tmp2103 = {tmp12[255]};
    assign tmp2104 = ~tmp2103;
    assign tmp2105 = tmp2102 ^ tmp2104;
    assign tmp2106 = {tmp2100[255]};
    assign tmp2107 = ~tmp2106;
    assign tmp2108 = tmp2105 ^ tmp2107;
    assign tmp2109 = {tmp13[255]};
    assign tmp2110 = {const_222_0};
    assign tmp2111 = {tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110, tmp2110};
    assign tmp2112 = {tmp2111, const_222_0};
    assign tmp2113 = tmp13 - tmp2112;
    assign tmp2114 = {tmp2113[256]};
    assign tmp2115 = {tmp13[255]};
    assign tmp2116 = ~tmp2115;
    assign tmp2117 = tmp2114 ^ tmp2116;
    assign tmp2118 = {tmp2112[255]};
    assign tmp2119 = ~tmp2118;
    assign tmp2120 = tmp2117 ^ tmp2119;
    assign tmp2121 = tmp2108 == tmp2120;
    assign tmp2122 = tmp2096 & tmp2121;
    assign tmp2123 = {tmp13[255]};
    assign tmp2124 = {const_223_0};
    assign tmp2125 = {tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124, tmp2124};
    assign tmp2126 = {tmp2125, const_223_0};
    assign tmp2127 = tmp13 - tmp2126;
    assign tmp2128 = {tmp2127[256]};
    assign tmp2129 = {tmp13[255]};
    assign tmp2130 = ~tmp2129;
    assign tmp2131 = tmp2128 ^ tmp2130;
    assign tmp2132 = {tmp2126[255]};
    assign tmp2133 = ~tmp2132;
    assign tmp2134 = tmp2131 ^ tmp2133;
    assign tmp2135 = {tmp14[255]};
    assign tmp2136 = {const_224_0};
    assign tmp2137 = {tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136, tmp2136};
    assign tmp2138 = {tmp2137, const_224_0};
    assign tmp2139 = tmp14 - tmp2138;
    assign tmp2140 = {tmp2139[256]};
    assign tmp2141 = {tmp14[255]};
    assign tmp2142 = ~tmp2141;
    assign tmp2143 = tmp2140 ^ tmp2142;
    assign tmp2144 = {tmp2138[255]};
    assign tmp2145 = ~tmp2144;
    assign tmp2146 = tmp2143 ^ tmp2145;
    assign tmp2147 = tmp2134 == tmp2146;
    assign tmp2148 = tmp2122 & tmp2147;
    assign tmp2149 = ~tmp35;
    assign tmp2150 = ~tmp36;
    assign tmp2151 = tmp2149 & tmp2150;
    assign tmp2152 = ~tmp57;
    assign tmp2153 = tmp2151 & tmp2152;
    assign tmp2154 = ~tmp1034;
    assign tmp2155 = tmp2153 & tmp2154;
    assign tmp2156 = tmp2155 & tmp2071;
    assign tmp2157 = {tmp15[255]};
    assign tmp2158 = {const_225_0};
    assign tmp2159 = {tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158, tmp2158};
    assign tmp2160 = {tmp2159, const_225_0};
    assign tmp2161 = tmp15 - tmp2160;
    assign tmp2162 = {tmp2161[256]};
    assign tmp2163 = {tmp15[255]};
    assign tmp2164 = ~tmp2163;
    assign tmp2165 = tmp2162 ^ tmp2164;
    assign tmp2166 = {tmp2160[255]};
    assign tmp2167 = ~tmp2166;
    assign tmp2168 = tmp2165 ^ tmp2167;
    assign tmp2169 = {tmp16[255]};
    assign tmp2170 = {const_226_0};
    assign tmp2171 = {tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170, tmp2170};
    assign tmp2172 = {tmp2171, const_226_0};
    assign tmp2173 = tmp16 - tmp2172;
    assign tmp2174 = {tmp2173[256]};
    assign tmp2175 = {tmp16[255]};
    assign tmp2176 = ~tmp2175;
    assign tmp2177 = tmp2174 ^ tmp2176;
    assign tmp2178 = {tmp2172[255]};
    assign tmp2179 = ~tmp2178;
    assign tmp2180 = tmp2177 ^ tmp2179;
    assign tmp2181 = tmp2168 == tmp2180;
    assign tmp2182 = {tmp16[255]};
    assign tmp2183 = {const_227_0};
    assign tmp2184 = {tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183, tmp2183};
    assign tmp2185 = {tmp2184, const_227_0};
    assign tmp2186 = tmp16 - tmp2185;
    assign tmp2187 = {tmp2186[256]};
    assign tmp2188 = {tmp16[255]};
    assign tmp2189 = ~tmp2188;
    assign tmp2190 = tmp2187 ^ tmp2189;
    assign tmp2191 = {tmp2185[255]};
    assign tmp2192 = ~tmp2191;
    assign tmp2193 = tmp2190 ^ tmp2192;
    assign tmp2194 = {tmp17[255]};
    assign tmp2195 = {const_228_0};
    assign tmp2196 = {tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195, tmp2195};
    assign tmp2197 = {tmp2196, const_228_0};
    assign tmp2198 = tmp17 - tmp2197;
    assign tmp2199 = {tmp2198[256]};
    assign tmp2200 = {tmp17[255]};
    assign tmp2201 = ~tmp2200;
    assign tmp2202 = tmp2199 ^ tmp2201;
    assign tmp2203 = {tmp2197[255]};
    assign tmp2204 = ~tmp2203;
    assign tmp2205 = tmp2202 ^ tmp2204;
    assign tmp2206 = tmp2193 == tmp2205;
    assign tmp2207 = tmp2181 & tmp2206;
    assign tmp2208 = {tmp17[255]};
    assign tmp2209 = {const_229_0};
    assign tmp2210 = {tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209, tmp2209};
    assign tmp2211 = {tmp2210, const_229_0};
    assign tmp2212 = tmp17 - tmp2211;
    assign tmp2213 = {tmp2212[256]};
    assign tmp2214 = {tmp17[255]};
    assign tmp2215 = ~tmp2214;
    assign tmp2216 = tmp2213 ^ tmp2215;
    assign tmp2217 = {tmp2211[255]};
    assign tmp2218 = ~tmp2217;
    assign tmp2219 = tmp2216 ^ tmp2218;
    assign tmp2220 = {tmp18[255]};
    assign tmp2221 = {const_230_0};
    assign tmp2222 = {tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221, tmp2221};
    assign tmp2223 = {tmp2222, const_230_0};
    assign tmp2224 = tmp18 - tmp2223;
    assign tmp2225 = {tmp2224[256]};
    assign tmp2226 = {tmp18[255]};
    assign tmp2227 = ~tmp2226;
    assign tmp2228 = tmp2225 ^ tmp2227;
    assign tmp2229 = {tmp2223[255]};
    assign tmp2230 = ~tmp2229;
    assign tmp2231 = tmp2228 ^ tmp2230;
    assign tmp2232 = tmp2219 == tmp2231;
    assign tmp2233 = tmp2207 & tmp2232;
    assign tmp2234 = ~tmp35;
    assign tmp2235 = ~tmp36;
    assign tmp2236 = tmp2234 & tmp2235;
    assign tmp2237 = ~tmp57;
    assign tmp2238 = tmp2236 & tmp2237;
    assign tmp2239 = ~tmp1034;
    assign tmp2240 = tmp2238 & tmp2239;
    assign tmp2241 = tmp2240 & tmp2071;
    assign tmp2242 = {const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0, const_232_0};
    assign tmp2243 = {tmp2242, const_231_0};
    assign tmp2244 = tmp15 == tmp2243;
    assign tmp2245 = {const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0, const_234_0};
    assign tmp2246 = {tmp2245, const_233_0};
    assign tmp2247 = tmp16 == tmp2246;
    assign tmp2248 = tmp2244 | tmp2247;
    assign tmp2249 = {const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0, const_236_0};
    assign tmp2250 = {tmp2249, const_235_0};
    assign tmp2251 = tmp17 == tmp2250;
    assign tmp2252 = tmp2248 | tmp2251;
    assign tmp2253 = {const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0, const_238_0};
    assign tmp2254 = {tmp2253, const_237_0};
    assign tmp2255 = tmp18 == tmp2254;
    assign tmp2256 = tmp2252 | tmp2255;
    assign tmp2257 = ~tmp35;
    assign tmp2258 = ~tmp36;
    assign tmp2259 = tmp2257 & tmp2258;
    assign tmp2260 = ~tmp57;
    assign tmp2261 = tmp2259 & tmp2260;
    assign tmp2262 = ~tmp1034;
    assign tmp2263 = tmp2261 & tmp2262;
    assign tmp2264 = tmp2263 & tmp2071;
    assign tmp2265 = tmp20 & tmp21;
    assign tmp2266 = ~tmp22;
    assign tmp2267 = tmp2265 & tmp2266;
    assign tmp2268 = ~tmp35;
    assign tmp2269 = ~tmp36;
    assign tmp2270 = tmp2268 & tmp2269;
    assign tmp2271 = ~tmp57;
    assign tmp2272 = tmp2270 & tmp2271;
    assign tmp2273 = ~tmp1034;
    assign tmp2274 = tmp2272 & tmp2273;
    assign tmp2275 = tmp2274 & tmp2071;
    assign tmp2276 = {tmp11[0]};
    assign tmp2277 = {tmp12[0]};
    assign tmp2278 = tmp2276 | tmp2277;
    assign tmp2279 = {tmp13[0]};
    assign tmp2280 = tmp2278 | tmp2279;
    assign tmp2281 = {tmp14[0]};
    assign tmp2282 = tmp2280 | tmp2281;
    assign tmp2283 = ~tmp2282;
    assign tmp2284 = ~tmp35;
    assign tmp2285 = ~tmp36;
    assign tmp2286 = tmp2284 & tmp2285;
    assign tmp2287 = ~tmp57;
    assign tmp2288 = tmp2286 & tmp2287;
    assign tmp2289 = ~tmp1034;
    assign tmp2290 = tmp2288 & tmp2289;
    assign tmp2291 = tmp2290 & tmp2071;
    assign tmp2292 = {tmp11[255]};
    assign tmp2293 = {const_239_0};
    assign tmp2294 = {tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293, tmp2293};
    assign tmp2295 = {tmp2294, const_239_0};
    assign tmp2296 = tmp11 - tmp2295;
    assign tmp2297 = {tmp2296[256]};
    assign tmp2298 = {tmp11[255]};
    assign tmp2299 = ~tmp2298;
    assign tmp2300 = tmp2297 ^ tmp2299;
    assign tmp2301 = {tmp2295[255]};
    assign tmp2302 = ~tmp2301;
    assign tmp2303 = tmp2300 ^ tmp2302;
    assign tmp2304 = tmp23 & tmp2303;
    assign tmp2305 = {tmp15[255]};
    assign tmp2306 = {const_240_0};
    assign tmp2307 = {tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306, tmp2306};
    assign tmp2308 = {tmp2307, const_240_0};
    assign tmp2309 = tmp15 - tmp2308;
    assign tmp2310 = {tmp2309[256]};
    assign tmp2311 = {tmp15[255]};
    assign tmp2312 = ~tmp2311;
    assign tmp2313 = tmp2310 ^ tmp2312;
    assign tmp2314 = {tmp2308[255]};
    assign tmp2315 = ~tmp2314;
    assign tmp2316 = tmp2313 ^ tmp2315;
    assign tmp2317 = tmp2304 & tmp2316;
    assign tmp2318 = tmp11 == _ver_out_tmp_83;
    assign tmp2319 = {const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0, const_243_0};
    assign tmp2320 = {tmp2319, const_242_0};
    assign tmp2321 = tmp2320 - tmp11;
    assign tmp2322 = {const_245_0, const_245_0};
    assign tmp2323 = {tmp2322, const_244_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp2324 = tmp2318 ? tmp2323 : tmp2321;
    assign tmp2325 = {tmp2324[255], tmp2324[254], tmp2324[253], tmp2324[252], tmp2324[251], tmp2324[250], tmp2324[249], tmp2324[248], tmp2324[247], tmp2324[246], tmp2324[245], tmp2324[244], tmp2324[243], tmp2324[242], tmp2324[241], tmp2324[240], tmp2324[239], tmp2324[238], tmp2324[237], tmp2324[236], tmp2324[235], tmp2324[234], tmp2324[233], tmp2324[232], tmp2324[231], tmp2324[230], tmp2324[229], tmp2324[228], tmp2324[227], tmp2324[226], tmp2324[225], tmp2324[224], tmp2324[223], tmp2324[222], tmp2324[221], tmp2324[220], tmp2324[219], tmp2324[218], tmp2324[217], tmp2324[216], tmp2324[215], tmp2324[214], tmp2324[213], tmp2324[212], tmp2324[211], tmp2324[210], tmp2324[209], tmp2324[208], tmp2324[207], tmp2324[206], tmp2324[205], tmp2324[204], tmp2324[203], tmp2324[202], tmp2324[201], tmp2324[200], tmp2324[199], tmp2324[198], tmp2324[197], tmp2324[196], tmp2324[195], tmp2324[194], tmp2324[193], tmp2324[192], tmp2324[191], tmp2324[190], tmp2324[189], tmp2324[188], tmp2324[187], tmp2324[186], tmp2324[185], tmp2324[184], tmp2324[183], tmp2324[182], tmp2324[181], tmp2324[180], tmp2324[179], tmp2324[178], tmp2324[177], tmp2324[176], tmp2324[175], tmp2324[174], tmp2324[173], tmp2324[172], tmp2324[171], tmp2324[170], tmp2324[169], tmp2324[168], tmp2324[167], tmp2324[166], tmp2324[165], tmp2324[164], tmp2324[163], tmp2324[162], tmp2324[161], tmp2324[160], tmp2324[159], tmp2324[158], tmp2324[157], tmp2324[156], tmp2324[155], tmp2324[154], tmp2324[153], tmp2324[152], tmp2324[151], tmp2324[150], tmp2324[149], tmp2324[148], tmp2324[147], tmp2324[146], tmp2324[145], tmp2324[144], tmp2324[143], tmp2324[142], tmp2324[141], tmp2324[140], tmp2324[139], tmp2324[138], tmp2324[137], tmp2324[136], tmp2324[135], tmp2324[134], tmp2324[133], tmp2324[132], tmp2324[131], tmp2324[130], tmp2324[129], tmp2324[128], tmp2324[127], tmp2324[126], tmp2324[125], tmp2324[124], tmp2324[123], tmp2324[122], tmp2324[121], tmp2324[120], tmp2324[119], tmp2324[118], tmp2324[117], tmp2324[116], tmp2324[115], tmp2324[114], tmp2324[113], tmp2324[112], tmp2324[111], tmp2324[110], tmp2324[109], tmp2324[108], tmp2324[107], tmp2324[106], tmp2324[105], tmp2324[104], tmp2324[103], tmp2324[102], tmp2324[101], tmp2324[100], tmp2324[99], tmp2324[98], tmp2324[97], tmp2324[96], tmp2324[95], tmp2324[94], tmp2324[93], tmp2324[92], tmp2324[91], tmp2324[90], tmp2324[89], tmp2324[88], tmp2324[87], tmp2324[86], tmp2324[85], tmp2324[84], tmp2324[83], tmp2324[82], tmp2324[81], tmp2324[80], tmp2324[79], tmp2324[78], tmp2324[77], tmp2324[76], tmp2324[75], tmp2324[74], tmp2324[73], tmp2324[72], tmp2324[71], tmp2324[70], tmp2324[69], tmp2324[68], tmp2324[67], tmp2324[66], tmp2324[65], tmp2324[64], tmp2324[63], tmp2324[62], tmp2324[61], tmp2324[60], tmp2324[59], tmp2324[58], tmp2324[57], tmp2324[56], tmp2324[55], tmp2324[54], tmp2324[53], tmp2324[52], tmp2324[51], tmp2324[50], tmp2324[49], tmp2324[48], tmp2324[47], tmp2324[46], tmp2324[45], tmp2324[44], tmp2324[43], tmp2324[42], tmp2324[41], tmp2324[40], tmp2324[39], tmp2324[38], tmp2324[37], tmp2324[36], tmp2324[35], tmp2324[34], tmp2324[33], tmp2324[32], tmp2324[31], tmp2324[30], tmp2324[29], tmp2324[28], tmp2324[27], tmp2324[26], tmp2324[25], tmp2324[24], tmp2324[23], tmp2324[22], tmp2324[21], tmp2324[20], tmp2324[19], tmp2324[18], tmp2324[17], tmp2324[16], tmp2324[15], tmp2324[14], tmp2324[13], tmp2324[12], tmp2324[11], tmp2324[10], tmp2324[9], tmp2324[8], tmp2324[7], tmp2324[6], tmp2324[5], tmp2324[4], tmp2324[3], tmp2324[2], tmp2324[1], tmp2324[0]};
    assign tmp2326 = ~tmp35;
    assign tmp2327 = ~tmp36;
    assign tmp2328 = tmp2326 & tmp2327;
    assign tmp2329 = ~tmp57;
    assign tmp2330 = tmp2328 & tmp2329;
    assign tmp2331 = ~tmp1034;
    assign tmp2332 = tmp2330 & tmp2331;
    assign tmp2333 = tmp2332 & tmp2071;
    assign tmp2334 = tmp2333 & tmp2317;
    assign tmp2335 = tmp12 == _ver_out_tmp_45;
    assign tmp2336 = {const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0, const_248_0};
    assign tmp2337 = {tmp2336, const_247_0};
    assign tmp2338 = tmp2337 - tmp12;
    assign tmp2339 = {const_250_0, const_250_0};
    assign tmp2340 = {tmp2339, const_249_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp2341 = tmp2335 ? tmp2340 : tmp2338;
    assign tmp2342 = {tmp2341[255], tmp2341[254], tmp2341[253], tmp2341[252], tmp2341[251], tmp2341[250], tmp2341[249], tmp2341[248], tmp2341[247], tmp2341[246], tmp2341[245], tmp2341[244], tmp2341[243], tmp2341[242], tmp2341[241], tmp2341[240], tmp2341[239], tmp2341[238], tmp2341[237], tmp2341[236], tmp2341[235], tmp2341[234], tmp2341[233], tmp2341[232], tmp2341[231], tmp2341[230], tmp2341[229], tmp2341[228], tmp2341[227], tmp2341[226], tmp2341[225], tmp2341[224], tmp2341[223], tmp2341[222], tmp2341[221], tmp2341[220], tmp2341[219], tmp2341[218], tmp2341[217], tmp2341[216], tmp2341[215], tmp2341[214], tmp2341[213], tmp2341[212], tmp2341[211], tmp2341[210], tmp2341[209], tmp2341[208], tmp2341[207], tmp2341[206], tmp2341[205], tmp2341[204], tmp2341[203], tmp2341[202], tmp2341[201], tmp2341[200], tmp2341[199], tmp2341[198], tmp2341[197], tmp2341[196], tmp2341[195], tmp2341[194], tmp2341[193], tmp2341[192], tmp2341[191], tmp2341[190], tmp2341[189], tmp2341[188], tmp2341[187], tmp2341[186], tmp2341[185], tmp2341[184], tmp2341[183], tmp2341[182], tmp2341[181], tmp2341[180], tmp2341[179], tmp2341[178], tmp2341[177], tmp2341[176], tmp2341[175], tmp2341[174], tmp2341[173], tmp2341[172], tmp2341[171], tmp2341[170], tmp2341[169], tmp2341[168], tmp2341[167], tmp2341[166], tmp2341[165], tmp2341[164], tmp2341[163], tmp2341[162], tmp2341[161], tmp2341[160], tmp2341[159], tmp2341[158], tmp2341[157], tmp2341[156], tmp2341[155], tmp2341[154], tmp2341[153], tmp2341[152], tmp2341[151], tmp2341[150], tmp2341[149], tmp2341[148], tmp2341[147], tmp2341[146], tmp2341[145], tmp2341[144], tmp2341[143], tmp2341[142], tmp2341[141], tmp2341[140], tmp2341[139], tmp2341[138], tmp2341[137], tmp2341[136], tmp2341[135], tmp2341[134], tmp2341[133], tmp2341[132], tmp2341[131], tmp2341[130], tmp2341[129], tmp2341[128], tmp2341[127], tmp2341[126], tmp2341[125], tmp2341[124], tmp2341[123], tmp2341[122], tmp2341[121], tmp2341[120], tmp2341[119], tmp2341[118], tmp2341[117], tmp2341[116], tmp2341[115], tmp2341[114], tmp2341[113], tmp2341[112], tmp2341[111], tmp2341[110], tmp2341[109], tmp2341[108], tmp2341[107], tmp2341[106], tmp2341[105], tmp2341[104], tmp2341[103], tmp2341[102], tmp2341[101], tmp2341[100], tmp2341[99], tmp2341[98], tmp2341[97], tmp2341[96], tmp2341[95], tmp2341[94], tmp2341[93], tmp2341[92], tmp2341[91], tmp2341[90], tmp2341[89], tmp2341[88], tmp2341[87], tmp2341[86], tmp2341[85], tmp2341[84], tmp2341[83], tmp2341[82], tmp2341[81], tmp2341[80], tmp2341[79], tmp2341[78], tmp2341[77], tmp2341[76], tmp2341[75], tmp2341[74], tmp2341[73], tmp2341[72], tmp2341[71], tmp2341[70], tmp2341[69], tmp2341[68], tmp2341[67], tmp2341[66], tmp2341[65], tmp2341[64], tmp2341[63], tmp2341[62], tmp2341[61], tmp2341[60], tmp2341[59], tmp2341[58], tmp2341[57], tmp2341[56], tmp2341[55], tmp2341[54], tmp2341[53], tmp2341[52], tmp2341[51], tmp2341[50], tmp2341[49], tmp2341[48], tmp2341[47], tmp2341[46], tmp2341[45], tmp2341[44], tmp2341[43], tmp2341[42], tmp2341[41], tmp2341[40], tmp2341[39], tmp2341[38], tmp2341[37], tmp2341[36], tmp2341[35], tmp2341[34], tmp2341[33], tmp2341[32], tmp2341[31], tmp2341[30], tmp2341[29], tmp2341[28], tmp2341[27], tmp2341[26], tmp2341[25], tmp2341[24], tmp2341[23], tmp2341[22], tmp2341[21], tmp2341[20], tmp2341[19], tmp2341[18], tmp2341[17], tmp2341[16], tmp2341[15], tmp2341[14], tmp2341[13], tmp2341[12], tmp2341[11], tmp2341[10], tmp2341[9], tmp2341[8], tmp2341[7], tmp2341[6], tmp2341[5], tmp2341[4], tmp2341[3], tmp2341[2], tmp2341[1], tmp2341[0]};
    assign tmp2343 = ~tmp35;
    assign tmp2344 = ~tmp36;
    assign tmp2345 = tmp2343 & tmp2344;
    assign tmp2346 = ~tmp57;
    assign tmp2347 = tmp2345 & tmp2346;
    assign tmp2348 = ~tmp1034;
    assign tmp2349 = tmp2347 & tmp2348;
    assign tmp2350 = tmp2349 & tmp2071;
    assign tmp2351 = tmp2350 & tmp2317;
    assign tmp2352 = tmp13 == _ver_out_tmp_86;
    assign tmp2353 = {const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0, const_253_0};
    assign tmp2354 = {tmp2353, const_252_0};
    assign tmp2355 = tmp2354 - tmp13;
    assign tmp2356 = {const_255_0, const_255_0};
    assign tmp2357 = {tmp2356, const_254_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp2358 = tmp2352 ? tmp2357 : tmp2355;
    assign tmp2359 = {tmp2358[255], tmp2358[254], tmp2358[253], tmp2358[252], tmp2358[251], tmp2358[250], tmp2358[249], tmp2358[248], tmp2358[247], tmp2358[246], tmp2358[245], tmp2358[244], tmp2358[243], tmp2358[242], tmp2358[241], tmp2358[240], tmp2358[239], tmp2358[238], tmp2358[237], tmp2358[236], tmp2358[235], tmp2358[234], tmp2358[233], tmp2358[232], tmp2358[231], tmp2358[230], tmp2358[229], tmp2358[228], tmp2358[227], tmp2358[226], tmp2358[225], tmp2358[224], tmp2358[223], tmp2358[222], tmp2358[221], tmp2358[220], tmp2358[219], tmp2358[218], tmp2358[217], tmp2358[216], tmp2358[215], tmp2358[214], tmp2358[213], tmp2358[212], tmp2358[211], tmp2358[210], tmp2358[209], tmp2358[208], tmp2358[207], tmp2358[206], tmp2358[205], tmp2358[204], tmp2358[203], tmp2358[202], tmp2358[201], tmp2358[200], tmp2358[199], tmp2358[198], tmp2358[197], tmp2358[196], tmp2358[195], tmp2358[194], tmp2358[193], tmp2358[192], tmp2358[191], tmp2358[190], tmp2358[189], tmp2358[188], tmp2358[187], tmp2358[186], tmp2358[185], tmp2358[184], tmp2358[183], tmp2358[182], tmp2358[181], tmp2358[180], tmp2358[179], tmp2358[178], tmp2358[177], tmp2358[176], tmp2358[175], tmp2358[174], tmp2358[173], tmp2358[172], tmp2358[171], tmp2358[170], tmp2358[169], tmp2358[168], tmp2358[167], tmp2358[166], tmp2358[165], tmp2358[164], tmp2358[163], tmp2358[162], tmp2358[161], tmp2358[160], tmp2358[159], tmp2358[158], tmp2358[157], tmp2358[156], tmp2358[155], tmp2358[154], tmp2358[153], tmp2358[152], tmp2358[151], tmp2358[150], tmp2358[149], tmp2358[148], tmp2358[147], tmp2358[146], tmp2358[145], tmp2358[144], tmp2358[143], tmp2358[142], tmp2358[141], tmp2358[140], tmp2358[139], tmp2358[138], tmp2358[137], tmp2358[136], tmp2358[135], tmp2358[134], tmp2358[133], tmp2358[132], tmp2358[131], tmp2358[130], tmp2358[129], tmp2358[128], tmp2358[127], tmp2358[126], tmp2358[125], tmp2358[124], tmp2358[123], tmp2358[122], tmp2358[121], tmp2358[120], tmp2358[119], tmp2358[118], tmp2358[117], tmp2358[116], tmp2358[115], tmp2358[114], tmp2358[113], tmp2358[112], tmp2358[111], tmp2358[110], tmp2358[109], tmp2358[108], tmp2358[107], tmp2358[106], tmp2358[105], tmp2358[104], tmp2358[103], tmp2358[102], tmp2358[101], tmp2358[100], tmp2358[99], tmp2358[98], tmp2358[97], tmp2358[96], tmp2358[95], tmp2358[94], tmp2358[93], tmp2358[92], tmp2358[91], tmp2358[90], tmp2358[89], tmp2358[88], tmp2358[87], tmp2358[86], tmp2358[85], tmp2358[84], tmp2358[83], tmp2358[82], tmp2358[81], tmp2358[80], tmp2358[79], tmp2358[78], tmp2358[77], tmp2358[76], tmp2358[75], tmp2358[74], tmp2358[73], tmp2358[72], tmp2358[71], tmp2358[70], tmp2358[69], tmp2358[68], tmp2358[67], tmp2358[66], tmp2358[65], tmp2358[64], tmp2358[63], tmp2358[62], tmp2358[61], tmp2358[60], tmp2358[59], tmp2358[58], tmp2358[57], tmp2358[56], tmp2358[55], tmp2358[54], tmp2358[53], tmp2358[52], tmp2358[51], tmp2358[50], tmp2358[49], tmp2358[48], tmp2358[47], tmp2358[46], tmp2358[45], tmp2358[44], tmp2358[43], tmp2358[42], tmp2358[41], tmp2358[40], tmp2358[39], tmp2358[38], tmp2358[37], tmp2358[36], tmp2358[35], tmp2358[34], tmp2358[33], tmp2358[32], tmp2358[31], tmp2358[30], tmp2358[29], tmp2358[28], tmp2358[27], tmp2358[26], tmp2358[25], tmp2358[24], tmp2358[23], tmp2358[22], tmp2358[21], tmp2358[20], tmp2358[19], tmp2358[18], tmp2358[17], tmp2358[16], tmp2358[15], tmp2358[14], tmp2358[13], tmp2358[12], tmp2358[11], tmp2358[10], tmp2358[9], tmp2358[8], tmp2358[7], tmp2358[6], tmp2358[5], tmp2358[4], tmp2358[3], tmp2358[2], tmp2358[1], tmp2358[0]};
    assign tmp2360 = ~tmp35;
    assign tmp2361 = ~tmp36;
    assign tmp2362 = tmp2360 & tmp2361;
    assign tmp2363 = ~tmp57;
    assign tmp2364 = tmp2362 & tmp2363;
    assign tmp2365 = ~tmp1034;
    assign tmp2366 = tmp2364 & tmp2365;
    assign tmp2367 = tmp2366 & tmp2071;
    assign tmp2368 = tmp2367 & tmp2317;
    assign tmp2369 = tmp14 == _ver_out_tmp_88;
    assign tmp2370 = {const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0, const_258_0};
    assign tmp2371 = {tmp2370, const_257_0};
    assign tmp2372 = tmp2371 - tmp14;
    assign tmp2373 = {const_260_0, const_260_0};
    assign tmp2374 = {tmp2373, const_259_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp2375 = tmp2369 ? tmp2374 : tmp2372;
    assign tmp2376 = {tmp2375[255], tmp2375[254], tmp2375[253], tmp2375[252], tmp2375[251], tmp2375[250], tmp2375[249], tmp2375[248], tmp2375[247], tmp2375[246], tmp2375[245], tmp2375[244], tmp2375[243], tmp2375[242], tmp2375[241], tmp2375[240], tmp2375[239], tmp2375[238], tmp2375[237], tmp2375[236], tmp2375[235], tmp2375[234], tmp2375[233], tmp2375[232], tmp2375[231], tmp2375[230], tmp2375[229], tmp2375[228], tmp2375[227], tmp2375[226], tmp2375[225], tmp2375[224], tmp2375[223], tmp2375[222], tmp2375[221], tmp2375[220], tmp2375[219], tmp2375[218], tmp2375[217], tmp2375[216], tmp2375[215], tmp2375[214], tmp2375[213], tmp2375[212], tmp2375[211], tmp2375[210], tmp2375[209], tmp2375[208], tmp2375[207], tmp2375[206], tmp2375[205], tmp2375[204], tmp2375[203], tmp2375[202], tmp2375[201], tmp2375[200], tmp2375[199], tmp2375[198], tmp2375[197], tmp2375[196], tmp2375[195], tmp2375[194], tmp2375[193], tmp2375[192], tmp2375[191], tmp2375[190], tmp2375[189], tmp2375[188], tmp2375[187], tmp2375[186], tmp2375[185], tmp2375[184], tmp2375[183], tmp2375[182], tmp2375[181], tmp2375[180], tmp2375[179], tmp2375[178], tmp2375[177], tmp2375[176], tmp2375[175], tmp2375[174], tmp2375[173], tmp2375[172], tmp2375[171], tmp2375[170], tmp2375[169], tmp2375[168], tmp2375[167], tmp2375[166], tmp2375[165], tmp2375[164], tmp2375[163], tmp2375[162], tmp2375[161], tmp2375[160], tmp2375[159], tmp2375[158], tmp2375[157], tmp2375[156], tmp2375[155], tmp2375[154], tmp2375[153], tmp2375[152], tmp2375[151], tmp2375[150], tmp2375[149], tmp2375[148], tmp2375[147], tmp2375[146], tmp2375[145], tmp2375[144], tmp2375[143], tmp2375[142], tmp2375[141], tmp2375[140], tmp2375[139], tmp2375[138], tmp2375[137], tmp2375[136], tmp2375[135], tmp2375[134], tmp2375[133], tmp2375[132], tmp2375[131], tmp2375[130], tmp2375[129], tmp2375[128], tmp2375[127], tmp2375[126], tmp2375[125], tmp2375[124], tmp2375[123], tmp2375[122], tmp2375[121], tmp2375[120], tmp2375[119], tmp2375[118], tmp2375[117], tmp2375[116], tmp2375[115], tmp2375[114], tmp2375[113], tmp2375[112], tmp2375[111], tmp2375[110], tmp2375[109], tmp2375[108], tmp2375[107], tmp2375[106], tmp2375[105], tmp2375[104], tmp2375[103], tmp2375[102], tmp2375[101], tmp2375[100], tmp2375[99], tmp2375[98], tmp2375[97], tmp2375[96], tmp2375[95], tmp2375[94], tmp2375[93], tmp2375[92], tmp2375[91], tmp2375[90], tmp2375[89], tmp2375[88], tmp2375[87], tmp2375[86], tmp2375[85], tmp2375[84], tmp2375[83], tmp2375[82], tmp2375[81], tmp2375[80], tmp2375[79], tmp2375[78], tmp2375[77], tmp2375[76], tmp2375[75], tmp2375[74], tmp2375[73], tmp2375[72], tmp2375[71], tmp2375[70], tmp2375[69], tmp2375[68], tmp2375[67], tmp2375[66], tmp2375[65], tmp2375[64], tmp2375[63], tmp2375[62], tmp2375[61], tmp2375[60], tmp2375[59], tmp2375[58], tmp2375[57], tmp2375[56], tmp2375[55], tmp2375[54], tmp2375[53], tmp2375[52], tmp2375[51], tmp2375[50], tmp2375[49], tmp2375[48], tmp2375[47], tmp2375[46], tmp2375[45], tmp2375[44], tmp2375[43], tmp2375[42], tmp2375[41], tmp2375[40], tmp2375[39], tmp2375[38], tmp2375[37], tmp2375[36], tmp2375[35], tmp2375[34], tmp2375[33], tmp2375[32], tmp2375[31], tmp2375[30], tmp2375[29], tmp2375[28], tmp2375[27], tmp2375[26], tmp2375[25], tmp2375[24], tmp2375[23], tmp2375[22], tmp2375[21], tmp2375[20], tmp2375[19], tmp2375[18], tmp2375[17], tmp2375[16], tmp2375[15], tmp2375[14], tmp2375[13], tmp2375[12], tmp2375[11], tmp2375[10], tmp2375[9], tmp2375[8], tmp2375[7], tmp2375[6], tmp2375[5], tmp2375[4], tmp2375[3], tmp2375[2], tmp2375[1], tmp2375[0]};
    assign tmp2377 = ~tmp35;
    assign tmp2378 = ~tmp36;
    assign tmp2379 = tmp2377 & tmp2378;
    assign tmp2380 = ~tmp57;
    assign tmp2381 = tmp2379 & tmp2380;
    assign tmp2382 = ~tmp1034;
    assign tmp2383 = tmp2381 & tmp2382;
    assign tmp2384 = tmp2383 & tmp2071;
    assign tmp2385 = tmp2384 & tmp2317;
    assign tmp2386 = tmp15 == _ver_out_tmp_89;
    assign tmp2387 = {const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0, const_263_0};
    assign tmp2388 = {tmp2387, const_262_0};
    assign tmp2389 = tmp2388 - tmp15;
    assign tmp2390 = {const_265_0, const_265_0};
    assign tmp2391 = {tmp2390, const_264_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp2392 = tmp2386 ? tmp2391 : tmp2389;
    assign tmp2393 = {tmp2392[255], tmp2392[254], tmp2392[253], tmp2392[252], tmp2392[251], tmp2392[250], tmp2392[249], tmp2392[248], tmp2392[247], tmp2392[246], tmp2392[245], tmp2392[244], tmp2392[243], tmp2392[242], tmp2392[241], tmp2392[240], tmp2392[239], tmp2392[238], tmp2392[237], tmp2392[236], tmp2392[235], tmp2392[234], tmp2392[233], tmp2392[232], tmp2392[231], tmp2392[230], tmp2392[229], tmp2392[228], tmp2392[227], tmp2392[226], tmp2392[225], tmp2392[224], tmp2392[223], tmp2392[222], tmp2392[221], tmp2392[220], tmp2392[219], tmp2392[218], tmp2392[217], tmp2392[216], tmp2392[215], tmp2392[214], tmp2392[213], tmp2392[212], tmp2392[211], tmp2392[210], tmp2392[209], tmp2392[208], tmp2392[207], tmp2392[206], tmp2392[205], tmp2392[204], tmp2392[203], tmp2392[202], tmp2392[201], tmp2392[200], tmp2392[199], tmp2392[198], tmp2392[197], tmp2392[196], tmp2392[195], tmp2392[194], tmp2392[193], tmp2392[192], tmp2392[191], tmp2392[190], tmp2392[189], tmp2392[188], tmp2392[187], tmp2392[186], tmp2392[185], tmp2392[184], tmp2392[183], tmp2392[182], tmp2392[181], tmp2392[180], tmp2392[179], tmp2392[178], tmp2392[177], tmp2392[176], tmp2392[175], tmp2392[174], tmp2392[173], tmp2392[172], tmp2392[171], tmp2392[170], tmp2392[169], tmp2392[168], tmp2392[167], tmp2392[166], tmp2392[165], tmp2392[164], tmp2392[163], tmp2392[162], tmp2392[161], tmp2392[160], tmp2392[159], tmp2392[158], tmp2392[157], tmp2392[156], tmp2392[155], tmp2392[154], tmp2392[153], tmp2392[152], tmp2392[151], tmp2392[150], tmp2392[149], tmp2392[148], tmp2392[147], tmp2392[146], tmp2392[145], tmp2392[144], tmp2392[143], tmp2392[142], tmp2392[141], tmp2392[140], tmp2392[139], tmp2392[138], tmp2392[137], tmp2392[136], tmp2392[135], tmp2392[134], tmp2392[133], tmp2392[132], tmp2392[131], tmp2392[130], tmp2392[129], tmp2392[128], tmp2392[127], tmp2392[126], tmp2392[125], tmp2392[124], tmp2392[123], tmp2392[122], tmp2392[121], tmp2392[120], tmp2392[119], tmp2392[118], tmp2392[117], tmp2392[116], tmp2392[115], tmp2392[114], tmp2392[113], tmp2392[112], tmp2392[111], tmp2392[110], tmp2392[109], tmp2392[108], tmp2392[107], tmp2392[106], tmp2392[105], tmp2392[104], tmp2392[103], tmp2392[102], tmp2392[101], tmp2392[100], tmp2392[99], tmp2392[98], tmp2392[97], tmp2392[96], tmp2392[95], tmp2392[94], tmp2392[93], tmp2392[92], tmp2392[91], tmp2392[90], tmp2392[89], tmp2392[88], tmp2392[87], tmp2392[86], tmp2392[85], tmp2392[84], tmp2392[83], tmp2392[82], tmp2392[81], tmp2392[80], tmp2392[79], tmp2392[78], tmp2392[77], tmp2392[76], tmp2392[75], tmp2392[74], tmp2392[73], tmp2392[72], tmp2392[71], tmp2392[70], tmp2392[69], tmp2392[68], tmp2392[67], tmp2392[66], tmp2392[65], tmp2392[64], tmp2392[63], tmp2392[62], tmp2392[61], tmp2392[60], tmp2392[59], tmp2392[58], tmp2392[57], tmp2392[56], tmp2392[55], tmp2392[54], tmp2392[53], tmp2392[52], tmp2392[51], tmp2392[50], tmp2392[49], tmp2392[48], tmp2392[47], tmp2392[46], tmp2392[45], tmp2392[44], tmp2392[43], tmp2392[42], tmp2392[41], tmp2392[40], tmp2392[39], tmp2392[38], tmp2392[37], tmp2392[36], tmp2392[35], tmp2392[34], tmp2392[33], tmp2392[32], tmp2392[31], tmp2392[30], tmp2392[29], tmp2392[28], tmp2392[27], tmp2392[26], tmp2392[25], tmp2392[24], tmp2392[23], tmp2392[22], tmp2392[21], tmp2392[20], tmp2392[19], tmp2392[18], tmp2392[17], tmp2392[16], tmp2392[15], tmp2392[14], tmp2392[13], tmp2392[12], tmp2392[11], tmp2392[10], tmp2392[9], tmp2392[8], tmp2392[7], tmp2392[6], tmp2392[5], tmp2392[4], tmp2392[3], tmp2392[2], tmp2392[1], tmp2392[0]};
    assign tmp2394 = ~tmp35;
    assign tmp2395 = ~tmp36;
    assign tmp2396 = tmp2394 & tmp2395;
    assign tmp2397 = ~tmp57;
    assign tmp2398 = tmp2396 & tmp2397;
    assign tmp2399 = ~tmp1034;
    assign tmp2400 = tmp2398 & tmp2399;
    assign tmp2401 = tmp2400 & tmp2071;
    assign tmp2402 = tmp2401 & tmp2317;
    assign tmp2403 = tmp16 == _ver_out_tmp_91;
    assign tmp2404 = {const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0, const_268_0};
    assign tmp2405 = {tmp2404, const_267_0};
    assign tmp2406 = tmp2405 - tmp16;
    assign tmp2407 = {const_270_0, const_270_0};
    assign tmp2408 = {tmp2407, const_269_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp2409 = tmp2403 ? tmp2408 : tmp2406;
    assign tmp2410 = {tmp2409[255], tmp2409[254], tmp2409[253], tmp2409[252], tmp2409[251], tmp2409[250], tmp2409[249], tmp2409[248], tmp2409[247], tmp2409[246], tmp2409[245], tmp2409[244], tmp2409[243], tmp2409[242], tmp2409[241], tmp2409[240], tmp2409[239], tmp2409[238], tmp2409[237], tmp2409[236], tmp2409[235], tmp2409[234], tmp2409[233], tmp2409[232], tmp2409[231], tmp2409[230], tmp2409[229], tmp2409[228], tmp2409[227], tmp2409[226], tmp2409[225], tmp2409[224], tmp2409[223], tmp2409[222], tmp2409[221], tmp2409[220], tmp2409[219], tmp2409[218], tmp2409[217], tmp2409[216], tmp2409[215], tmp2409[214], tmp2409[213], tmp2409[212], tmp2409[211], tmp2409[210], tmp2409[209], tmp2409[208], tmp2409[207], tmp2409[206], tmp2409[205], tmp2409[204], tmp2409[203], tmp2409[202], tmp2409[201], tmp2409[200], tmp2409[199], tmp2409[198], tmp2409[197], tmp2409[196], tmp2409[195], tmp2409[194], tmp2409[193], tmp2409[192], tmp2409[191], tmp2409[190], tmp2409[189], tmp2409[188], tmp2409[187], tmp2409[186], tmp2409[185], tmp2409[184], tmp2409[183], tmp2409[182], tmp2409[181], tmp2409[180], tmp2409[179], tmp2409[178], tmp2409[177], tmp2409[176], tmp2409[175], tmp2409[174], tmp2409[173], tmp2409[172], tmp2409[171], tmp2409[170], tmp2409[169], tmp2409[168], tmp2409[167], tmp2409[166], tmp2409[165], tmp2409[164], tmp2409[163], tmp2409[162], tmp2409[161], tmp2409[160], tmp2409[159], tmp2409[158], tmp2409[157], tmp2409[156], tmp2409[155], tmp2409[154], tmp2409[153], tmp2409[152], tmp2409[151], tmp2409[150], tmp2409[149], tmp2409[148], tmp2409[147], tmp2409[146], tmp2409[145], tmp2409[144], tmp2409[143], tmp2409[142], tmp2409[141], tmp2409[140], tmp2409[139], tmp2409[138], tmp2409[137], tmp2409[136], tmp2409[135], tmp2409[134], tmp2409[133], tmp2409[132], tmp2409[131], tmp2409[130], tmp2409[129], tmp2409[128], tmp2409[127], tmp2409[126], tmp2409[125], tmp2409[124], tmp2409[123], tmp2409[122], tmp2409[121], tmp2409[120], tmp2409[119], tmp2409[118], tmp2409[117], tmp2409[116], tmp2409[115], tmp2409[114], tmp2409[113], tmp2409[112], tmp2409[111], tmp2409[110], tmp2409[109], tmp2409[108], tmp2409[107], tmp2409[106], tmp2409[105], tmp2409[104], tmp2409[103], tmp2409[102], tmp2409[101], tmp2409[100], tmp2409[99], tmp2409[98], tmp2409[97], tmp2409[96], tmp2409[95], tmp2409[94], tmp2409[93], tmp2409[92], tmp2409[91], tmp2409[90], tmp2409[89], tmp2409[88], tmp2409[87], tmp2409[86], tmp2409[85], tmp2409[84], tmp2409[83], tmp2409[82], tmp2409[81], tmp2409[80], tmp2409[79], tmp2409[78], tmp2409[77], tmp2409[76], tmp2409[75], tmp2409[74], tmp2409[73], tmp2409[72], tmp2409[71], tmp2409[70], tmp2409[69], tmp2409[68], tmp2409[67], tmp2409[66], tmp2409[65], tmp2409[64], tmp2409[63], tmp2409[62], tmp2409[61], tmp2409[60], tmp2409[59], tmp2409[58], tmp2409[57], tmp2409[56], tmp2409[55], tmp2409[54], tmp2409[53], tmp2409[52], tmp2409[51], tmp2409[50], tmp2409[49], tmp2409[48], tmp2409[47], tmp2409[46], tmp2409[45], tmp2409[44], tmp2409[43], tmp2409[42], tmp2409[41], tmp2409[40], tmp2409[39], tmp2409[38], tmp2409[37], tmp2409[36], tmp2409[35], tmp2409[34], tmp2409[33], tmp2409[32], tmp2409[31], tmp2409[30], tmp2409[29], tmp2409[28], tmp2409[27], tmp2409[26], tmp2409[25], tmp2409[24], tmp2409[23], tmp2409[22], tmp2409[21], tmp2409[20], tmp2409[19], tmp2409[18], tmp2409[17], tmp2409[16], tmp2409[15], tmp2409[14], tmp2409[13], tmp2409[12], tmp2409[11], tmp2409[10], tmp2409[9], tmp2409[8], tmp2409[7], tmp2409[6], tmp2409[5], tmp2409[4], tmp2409[3], tmp2409[2], tmp2409[1], tmp2409[0]};
    assign tmp2411 = ~tmp35;
    assign tmp2412 = ~tmp36;
    assign tmp2413 = tmp2411 & tmp2412;
    assign tmp2414 = ~tmp57;
    assign tmp2415 = tmp2413 & tmp2414;
    assign tmp2416 = ~tmp1034;
    assign tmp2417 = tmp2415 & tmp2416;
    assign tmp2418 = tmp2417 & tmp2071;
    assign tmp2419 = tmp2418 & tmp2317;
    assign tmp2420 = tmp17 == _ver_out_tmp_80;
    assign tmp2421 = {const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0, const_273_0};
    assign tmp2422 = {tmp2421, const_272_0};
    assign tmp2423 = tmp2422 - tmp17;
    assign tmp2424 = {const_275_0, const_275_0};
    assign tmp2425 = {tmp2424, const_274_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp2426 = tmp2420 ? tmp2425 : tmp2423;
    assign tmp2427 = {tmp2426[255], tmp2426[254], tmp2426[253], tmp2426[252], tmp2426[251], tmp2426[250], tmp2426[249], tmp2426[248], tmp2426[247], tmp2426[246], tmp2426[245], tmp2426[244], tmp2426[243], tmp2426[242], tmp2426[241], tmp2426[240], tmp2426[239], tmp2426[238], tmp2426[237], tmp2426[236], tmp2426[235], tmp2426[234], tmp2426[233], tmp2426[232], tmp2426[231], tmp2426[230], tmp2426[229], tmp2426[228], tmp2426[227], tmp2426[226], tmp2426[225], tmp2426[224], tmp2426[223], tmp2426[222], tmp2426[221], tmp2426[220], tmp2426[219], tmp2426[218], tmp2426[217], tmp2426[216], tmp2426[215], tmp2426[214], tmp2426[213], tmp2426[212], tmp2426[211], tmp2426[210], tmp2426[209], tmp2426[208], tmp2426[207], tmp2426[206], tmp2426[205], tmp2426[204], tmp2426[203], tmp2426[202], tmp2426[201], tmp2426[200], tmp2426[199], tmp2426[198], tmp2426[197], tmp2426[196], tmp2426[195], tmp2426[194], tmp2426[193], tmp2426[192], tmp2426[191], tmp2426[190], tmp2426[189], tmp2426[188], tmp2426[187], tmp2426[186], tmp2426[185], tmp2426[184], tmp2426[183], tmp2426[182], tmp2426[181], tmp2426[180], tmp2426[179], tmp2426[178], tmp2426[177], tmp2426[176], tmp2426[175], tmp2426[174], tmp2426[173], tmp2426[172], tmp2426[171], tmp2426[170], tmp2426[169], tmp2426[168], tmp2426[167], tmp2426[166], tmp2426[165], tmp2426[164], tmp2426[163], tmp2426[162], tmp2426[161], tmp2426[160], tmp2426[159], tmp2426[158], tmp2426[157], tmp2426[156], tmp2426[155], tmp2426[154], tmp2426[153], tmp2426[152], tmp2426[151], tmp2426[150], tmp2426[149], tmp2426[148], tmp2426[147], tmp2426[146], tmp2426[145], tmp2426[144], tmp2426[143], tmp2426[142], tmp2426[141], tmp2426[140], tmp2426[139], tmp2426[138], tmp2426[137], tmp2426[136], tmp2426[135], tmp2426[134], tmp2426[133], tmp2426[132], tmp2426[131], tmp2426[130], tmp2426[129], tmp2426[128], tmp2426[127], tmp2426[126], tmp2426[125], tmp2426[124], tmp2426[123], tmp2426[122], tmp2426[121], tmp2426[120], tmp2426[119], tmp2426[118], tmp2426[117], tmp2426[116], tmp2426[115], tmp2426[114], tmp2426[113], tmp2426[112], tmp2426[111], tmp2426[110], tmp2426[109], tmp2426[108], tmp2426[107], tmp2426[106], tmp2426[105], tmp2426[104], tmp2426[103], tmp2426[102], tmp2426[101], tmp2426[100], tmp2426[99], tmp2426[98], tmp2426[97], tmp2426[96], tmp2426[95], tmp2426[94], tmp2426[93], tmp2426[92], tmp2426[91], tmp2426[90], tmp2426[89], tmp2426[88], tmp2426[87], tmp2426[86], tmp2426[85], tmp2426[84], tmp2426[83], tmp2426[82], tmp2426[81], tmp2426[80], tmp2426[79], tmp2426[78], tmp2426[77], tmp2426[76], tmp2426[75], tmp2426[74], tmp2426[73], tmp2426[72], tmp2426[71], tmp2426[70], tmp2426[69], tmp2426[68], tmp2426[67], tmp2426[66], tmp2426[65], tmp2426[64], tmp2426[63], tmp2426[62], tmp2426[61], tmp2426[60], tmp2426[59], tmp2426[58], tmp2426[57], tmp2426[56], tmp2426[55], tmp2426[54], tmp2426[53], tmp2426[52], tmp2426[51], tmp2426[50], tmp2426[49], tmp2426[48], tmp2426[47], tmp2426[46], tmp2426[45], tmp2426[44], tmp2426[43], tmp2426[42], tmp2426[41], tmp2426[40], tmp2426[39], tmp2426[38], tmp2426[37], tmp2426[36], tmp2426[35], tmp2426[34], tmp2426[33], tmp2426[32], tmp2426[31], tmp2426[30], tmp2426[29], tmp2426[28], tmp2426[27], tmp2426[26], tmp2426[25], tmp2426[24], tmp2426[23], tmp2426[22], tmp2426[21], tmp2426[20], tmp2426[19], tmp2426[18], tmp2426[17], tmp2426[16], tmp2426[15], tmp2426[14], tmp2426[13], tmp2426[12], tmp2426[11], tmp2426[10], tmp2426[9], tmp2426[8], tmp2426[7], tmp2426[6], tmp2426[5], tmp2426[4], tmp2426[3], tmp2426[2], tmp2426[1], tmp2426[0]};
    assign tmp2428 = ~tmp35;
    assign tmp2429 = ~tmp36;
    assign tmp2430 = tmp2428 & tmp2429;
    assign tmp2431 = ~tmp57;
    assign tmp2432 = tmp2430 & tmp2431;
    assign tmp2433 = ~tmp1034;
    assign tmp2434 = tmp2432 & tmp2433;
    assign tmp2435 = tmp2434 & tmp2071;
    assign tmp2436 = tmp2435 & tmp2317;
    assign tmp2437 = tmp18 == _ver_out_tmp_59;
    assign tmp2438 = {const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0, const_278_0};
    assign tmp2439 = {tmp2438, const_277_0};
    assign tmp2440 = tmp2439 - tmp18;
    assign tmp2441 = {const_280_0, const_280_0};
    assign tmp2442 = {tmp2441, const_279_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp2443 = tmp2437 ? tmp2442 : tmp2440;
    assign tmp2444 = {tmp2443[255], tmp2443[254], tmp2443[253], tmp2443[252], tmp2443[251], tmp2443[250], tmp2443[249], tmp2443[248], tmp2443[247], tmp2443[246], tmp2443[245], tmp2443[244], tmp2443[243], tmp2443[242], tmp2443[241], tmp2443[240], tmp2443[239], tmp2443[238], tmp2443[237], tmp2443[236], tmp2443[235], tmp2443[234], tmp2443[233], tmp2443[232], tmp2443[231], tmp2443[230], tmp2443[229], tmp2443[228], tmp2443[227], tmp2443[226], tmp2443[225], tmp2443[224], tmp2443[223], tmp2443[222], tmp2443[221], tmp2443[220], tmp2443[219], tmp2443[218], tmp2443[217], tmp2443[216], tmp2443[215], tmp2443[214], tmp2443[213], tmp2443[212], tmp2443[211], tmp2443[210], tmp2443[209], tmp2443[208], tmp2443[207], tmp2443[206], tmp2443[205], tmp2443[204], tmp2443[203], tmp2443[202], tmp2443[201], tmp2443[200], tmp2443[199], tmp2443[198], tmp2443[197], tmp2443[196], tmp2443[195], tmp2443[194], tmp2443[193], tmp2443[192], tmp2443[191], tmp2443[190], tmp2443[189], tmp2443[188], tmp2443[187], tmp2443[186], tmp2443[185], tmp2443[184], tmp2443[183], tmp2443[182], tmp2443[181], tmp2443[180], tmp2443[179], tmp2443[178], tmp2443[177], tmp2443[176], tmp2443[175], tmp2443[174], tmp2443[173], tmp2443[172], tmp2443[171], tmp2443[170], tmp2443[169], tmp2443[168], tmp2443[167], tmp2443[166], tmp2443[165], tmp2443[164], tmp2443[163], tmp2443[162], tmp2443[161], tmp2443[160], tmp2443[159], tmp2443[158], tmp2443[157], tmp2443[156], tmp2443[155], tmp2443[154], tmp2443[153], tmp2443[152], tmp2443[151], tmp2443[150], tmp2443[149], tmp2443[148], tmp2443[147], tmp2443[146], tmp2443[145], tmp2443[144], tmp2443[143], tmp2443[142], tmp2443[141], tmp2443[140], tmp2443[139], tmp2443[138], tmp2443[137], tmp2443[136], tmp2443[135], tmp2443[134], tmp2443[133], tmp2443[132], tmp2443[131], tmp2443[130], tmp2443[129], tmp2443[128], tmp2443[127], tmp2443[126], tmp2443[125], tmp2443[124], tmp2443[123], tmp2443[122], tmp2443[121], tmp2443[120], tmp2443[119], tmp2443[118], tmp2443[117], tmp2443[116], tmp2443[115], tmp2443[114], tmp2443[113], tmp2443[112], tmp2443[111], tmp2443[110], tmp2443[109], tmp2443[108], tmp2443[107], tmp2443[106], tmp2443[105], tmp2443[104], tmp2443[103], tmp2443[102], tmp2443[101], tmp2443[100], tmp2443[99], tmp2443[98], tmp2443[97], tmp2443[96], tmp2443[95], tmp2443[94], tmp2443[93], tmp2443[92], tmp2443[91], tmp2443[90], tmp2443[89], tmp2443[88], tmp2443[87], tmp2443[86], tmp2443[85], tmp2443[84], tmp2443[83], tmp2443[82], tmp2443[81], tmp2443[80], tmp2443[79], tmp2443[78], tmp2443[77], tmp2443[76], tmp2443[75], tmp2443[74], tmp2443[73], tmp2443[72], tmp2443[71], tmp2443[70], tmp2443[69], tmp2443[68], tmp2443[67], tmp2443[66], tmp2443[65], tmp2443[64], tmp2443[63], tmp2443[62], tmp2443[61], tmp2443[60], tmp2443[59], tmp2443[58], tmp2443[57], tmp2443[56], tmp2443[55], tmp2443[54], tmp2443[53], tmp2443[52], tmp2443[51], tmp2443[50], tmp2443[49], tmp2443[48], tmp2443[47], tmp2443[46], tmp2443[45], tmp2443[44], tmp2443[43], tmp2443[42], tmp2443[41], tmp2443[40], tmp2443[39], tmp2443[38], tmp2443[37], tmp2443[36], tmp2443[35], tmp2443[34], tmp2443[33], tmp2443[32], tmp2443[31], tmp2443[30], tmp2443[29], tmp2443[28], tmp2443[27], tmp2443[26], tmp2443[25], tmp2443[24], tmp2443[23], tmp2443[22], tmp2443[21], tmp2443[20], tmp2443[19], tmp2443[18], tmp2443[17], tmp2443[16], tmp2443[15], tmp2443[14], tmp2443[13], tmp2443[12], tmp2443[11], tmp2443[10], tmp2443[9], tmp2443[8], tmp2443[7], tmp2443[6], tmp2443[5], tmp2443[4], tmp2443[3], tmp2443[2], tmp2443[1], tmp2443[0]};
    assign tmp2445 = ~tmp35;
    assign tmp2446 = ~tmp36;
    assign tmp2447 = tmp2445 & tmp2446;
    assign tmp2448 = ~tmp57;
    assign tmp2449 = tmp2447 & tmp2448;
    assign tmp2450 = ~tmp1034;
    assign tmp2451 = tmp2449 & tmp2450;
    assign tmp2452 = tmp2451 & tmp2071;
    assign tmp2453 = tmp2452 & tmp2317;
    assign tmp2454 = {tmp11[255]};
    assign tmp2455 = {const_281_0};
    assign tmp2456 = {tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455, tmp2455};
    assign tmp2457 = {tmp2456, const_281_0};
    assign tmp2458 = tmp11 - tmp2457;
    assign tmp2459 = {tmp2458[256]};
    assign tmp2460 = {tmp11[255]};
    assign tmp2461 = ~tmp2460;
    assign tmp2462 = tmp2459 ^ tmp2461;
    assign tmp2463 = {tmp2457[255]};
    assign tmp2464 = ~tmp2463;
    assign tmp2465 = tmp2462 ^ tmp2464;
    assign tmp2466 = {tmp15[255]};
    assign tmp2467 = {const_282_0};
    assign tmp2468 = {tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467, tmp2467};
    assign tmp2469 = {tmp2468, const_282_0};
    assign tmp2470 = tmp15 - tmp2469;
    assign tmp2471 = {tmp2470[256]};
    assign tmp2472 = {tmp15[255]};
    assign tmp2473 = ~tmp2472;
    assign tmp2474 = tmp2471 ^ tmp2473;
    assign tmp2475 = {tmp2469[255]};
    assign tmp2476 = ~tmp2475;
    assign tmp2477 = tmp2474 ^ tmp2476;
    assign tmp2478 = tmp2465 & tmp2477;
    assign tmp2479 = ~tmp2478;
    assign tmp2480 = tmp23 & tmp2479;
    assign tmp2481 = ~tmp35;
    assign tmp2482 = ~tmp36;
    assign tmp2483 = tmp2481 & tmp2482;
    assign tmp2484 = ~tmp57;
    assign tmp2485 = tmp2483 & tmp2484;
    assign tmp2486 = ~tmp1034;
    assign tmp2487 = tmp2485 & tmp2486;
    assign tmp2488 = tmp2487 & tmp2071;
    assign tmp2489 = ~tmp2317;
    assign tmp2490 = tmp2488 & tmp2489;
    assign tmp2491 = tmp2490 & tmp2480;
    assign tmp2492 = ~tmp35;
    assign tmp2493 = ~tmp36;
    assign tmp2494 = tmp2492 & tmp2493;
    assign tmp2495 = ~tmp57;
    assign tmp2496 = tmp2494 & tmp2495;
    assign tmp2497 = ~tmp1034;
    assign tmp2498 = tmp2496 & tmp2497;
    assign tmp2499 = tmp2498 & tmp2071;
    assign tmp2500 = ~tmp2317;
    assign tmp2501 = tmp2499 & tmp2500;
    assign tmp2502 = tmp2501 & tmp2480;
    assign tmp2503 = ~tmp35;
    assign tmp2504 = ~tmp36;
    assign tmp2505 = tmp2503 & tmp2504;
    assign tmp2506 = ~tmp57;
    assign tmp2507 = tmp2505 & tmp2506;
    assign tmp2508 = ~tmp1034;
    assign tmp2509 = tmp2507 & tmp2508;
    assign tmp2510 = tmp2509 & tmp2071;
    assign tmp2511 = ~tmp2317;
    assign tmp2512 = tmp2510 & tmp2511;
    assign tmp2513 = tmp2512 & tmp2480;
    assign tmp2514 = ~tmp35;
    assign tmp2515 = ~tmp36;
    assign tmp2516 = tmp2514 & tmp2515;
    assign tmp2517 = ~tmp57;
    assign tmp2518 = tmp2516 & tmp2517;
    assign tmp2519 = ~tmp1034;
    assign tmp2520 = tmp2518 & tmp2519;
    assign tmp2521 = tmp2520 & tmp2071;
    assign tmp2522 = ~tmp2317;
    assign tmp2523 = tmp2521 & tmp2522;
    assign tmp2524 = tmp2523 & tmp2480;
    assign tmp2525 = ~tmp35;
    assign tmp2526 = ~tmp36;
    assign tmp2527 = tmp2525 & tmp2526;
    assign tmp2528 = ~tmp57;
    assign tmp2529 = tmp2527 & tmp2528;
    assign tmp2530 = ~tmp1034;
    assign tmp2531 = tmp2529 & tmp2530;
    assign tmp2532 = tmp2531 & tmp2071;
    assign tmp2533 = ~tmp2317;
    assign tmp2534 = tmp2532 & tmp2533;
    assign tmp2535 = tmp2534 & tmp2480;
    assign tmp2536 = ~tmp35;
    assign tmp2537 = ~tmp36;
    assign tmp2538 = tmp2536 & tmp2537;
    assign tmp2539 = ~tmp57;
    assign tmp2540 = tmp2538 & tmp2539;
    assign tmp2541 = ~tmp1034;
    assign tmp2542 = tmp2540 & tmp2541;
    assign tmp2543 = tmp2542 & tmp2071;
    assign tmp2544 = ~tmp2317;
    assign tmp2545 = tmp2543 & tmp2544;
    assign tmp2546 = tmp2545 & tmp2480;
    assign tmp2547 = ~tmp35;
    assign tmp2548 = ~tmp36;
    assign tmp2549 = tmp2547 & tmp2548;
    assign tmp2550 = ~tmp57;
    assign tmp2551 = tmp2549 & tmp2550;
    assign tmp2552 = ~tmp1034;
    assign tmp2553 = tmp2551 & tmp2552;
    assign tmp2554 = tmp2553 & tmp2071;
    assign tmp2555 = ~tmp2317;
    assign tmp2556 = tmp2554 & tmp2555;
    assign tmp2557 = tmp2556 & tmp2480;
    assign tmp2558 = ~tmp35;
    assign tmp2559 = ~tmp36;
    assign tmp2560 = tmp2558 & tmp2559;
    assign tmp2561 = ~tmp57;
    assign tmp2562 = tmp2560 & tmp2561;
    assign tmp2563 = ~tmp1034;
    assign tmp2564 = tmp2562 & tmp2563;
    assign tmp2565 = tmp2564 & tmp2071;
    assign tmp2566 = ~tmp2317;
    assign tmp2567 = tmp2565 & tmp2566;
    assign tmp2568 = tmp2567 & tmp2480;
    assign tmp2569 = {const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0, const_284_0};
    assign tmp2570 = {tmp2569, const_283_0};
    assign tmp2571 = tmp15 == tmp2570;
    assign tmp2572 = {const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0, const_286_0};
    assign tmp2573 = {tmp2572, const_285_0};
    assign tmp2574 = tmp16 == tmp2573;
    assign tmp2575 = tmp2571 & tmp2574;
    assign tmp2576 = {const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0, const_288_0};
    assign tmp2577 = {tmp2576, const_287_0};
    assign tmp2578 = tmp17 == tmp2577;
    assign tmp2579 = tmp2575 & tmp2578;
    assign tmp2580 = {const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0, const_290_0};
    assign tmp2581 = {tmp2580, const_289_0};
    assign tmp2582 = tmp18 == tmp2581;
    assign tmp2583 = tmp2579 & tmp2582;
    assign tmp2584 = ~tmp35;
    assign tmp2585 = ~tmp36;
    assign tmp2586 = tmp2584 & tmp2585;
    assign tmp2587 = ~tmp57;
    assign tmp2588 = tmp2586 & tmp2587;
    assign tmp2589 = ~tmp1034;
    assign tmp2590 = tmp2588 & tmp2589;
    assign tmp2591 = tmp2590 & tmp2071;
    assign tmp2592 = tmp2591 & tmp2583;
    assign tmp2593 = ~tmp35;
    assign tmp2594 = ~tmp36;
    assign tmp2595 = tmp2593 & tmp2594;
    assign tmp2596 = ~tmp57;
    assign tmp2597 = tmp2595 & tmp2596;
    assign tmp2598 = ~tmp1034;
    assign tmp2599 = tmp2597 & tmp2598;
    assign tmp2600 = tmp2599 & tmp2071;
    assign tmp2601 = tmp2600 & tmp2583;
    assign tmp2602 = {tmp11[255]};
    assign tmp2603 = {const_293_0};
    assign tmp2604 = {tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603, tmp2603};
    assign tmp2605 = {tmp2604, const_293_0};
    assign tmp2606 = tmp11 - tmp2605;
    assign tmp2607 = {tmp2606[256]};
    assign tmp2608 = {tmp11[255]};
    assign tmp2609 = ~tmp2608;
    assign tmp2610 = tmp2607 ^ tmp2609;
    assign tmp2611 = {tmp2605[255]};
    assign tmp2612 = ~tmp2611;
    assign tmp2613 = tmp2610 ^ tmp2612;
    assign tmp2614 = {tmp15[255]};
    assign tmp2615 = {const_294_0};
    assign tmp2616 = {tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615, tmp2615};
    assign tmp2617 = {tmp2616, const_294_0};
    assign tmp2618 = tmp15 - tmp2617;
    assign tmp2619 = {tmp2618[256]};
    assign tmp2620 = {tmp15[255]};
    assign tmp2621 = ~tmp2620;
    assign tmp2622 = tmp2619 ^ tmp2621;
    assign tmp2623 = {tmp2617[255]};
    assign tmp2624 = ~tmp2623;
    assign tmp2625 = tmp2622 ^ tmp2624;
    assign tmp2626 = tmp2613 == tmp2625;
    assign tmp2627 = ~tmp2626;
    assign tmp2628 = ~tmp35;
    assign tmp2629 = ~tmp36;
    assign tmp2630 = tmp2628 & tmp2629;
    assign tmp2631 = ~tmp57;
    assign tmp2632 = tmp2630 & tmp2631;
    assign tmp2633 = ~tmp1034;
    assign tmp2634 = tmp2632 & tmp2633;
    assign tmp2635 = tmp2634 & tmp2071;
    assign tmp2636 = ~tmp2583;
    assign tmp2637 = tmp2635 & tmp2636;
    assign tmp2638 = tmp2637 & tmp23;
    assign tmp2639 = tmp2638 & tmp2627;
    assign tmp2640 = ~tmp35;
    assign tmp2641 = ~tmp36;
    assign tmp2642 = tmp2640 & tmp2641;
    assign tmp2643 = ~tmp57;
    assign tmp2644 = tmp2642 & tmp2643;
    assign tmp2645 = ~tmp1034;
    assign tmp2646 = tmp2644 & tmp2645;
    assign tmp2647 = tmp2646 & tmp2071;
    assign tmp2648 = ~tmp2583;
    assign tmp2649 = tmp2647 & tmp2648;
    assign tmp2650 = tmp2649 & tmp23;
    assign tmp2651 = tmp2650 & tmp2627;
    assign tmp2652 = tmp11 == _ver_out_tmp_63;
    assign tmp2653 = {const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0, const_299_0};
    assign tmp2654 = {tmp2653, const_298_0};
    assign tmp2655 = tmp2654 - tmp11;
    assign tmp2656 = {const_301_0, const_301_0};
    assign tmp2657 = {tmp2656, const_300_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp2658 = tmp2652 ? tmp2657 : tmp2655;
    assign tmp2659 = {tmp2658[255], tmp2658[254], tmp2658[253], tmp2658[252], tmp2658[251], tmp2658[250], tmp2658[249], tmp2658[248], tmp2658[247], tmp2658[246], tmp2658[245], tmp2658[244], tmp2658[243], tmp2658[242], tmp2658[241], tmp2658[240], tmp2658[239], tmp2658[238], tmp2658[237], tmp2658[236], tmp2658[235], tmp2658[234], tmp2658[233], tmp2658[232], tmp2658[231], tmp2658[230], tmp2658[229], tmp2658[228], tmp2658[227], tmp2658[226], tmp2658[225], tmp2658[224], tmp2658[223], tmp2658[222], tmp2658[221], tmp2658[220], tmp2658[219], tmp2658[218], tmp2658[217], tmp2658[216], tmp2658[215], tmp2658[214], tmp2658[213], tmp2658[212], tmp2658[211], tmp2658[210], tmp2658[209], tmp2658[208], tmp2658[207], tmp2658[206], tmp2658[205], tmp2658[204], tmp2658[203], tmp2658[202], tmp2658[201], tmp2658[200], tmp2658[199], tmp2658[198], tmp2658[197], tmp2658[196], tmp2658[195], tmp2658[194], tmp2658[193], tmp2658[192], tmp2658[191], tmp2658[190], tmp2658[189], tmp2658[188], tmp2658[187], tmp2658[186], tmp2658[185], tmp2658[184], tmp2658[183], tmp2658[182], tmp2658[181], tmp2658[180], tmp2658[179], tmp2658[178], tmp2658[177], tmp2658[176], tmp2658[175], tmp2658[174], tmp2658[173], tmp2658[172], tmp2658[171], tmp2658[170], tmp2658[169], tmp2658[168], tmp2658[167], tmp2658[166], tmp2658[165], tmp2658[164], tmp2658[163], tmp2658[162], tmp2658[161], tmp2658[160], tmp2658[159], tmp2658[158], tmp2658[157], tmp2658[156], tmp2658[155], tmp2658[154], tmp2658[153], tmp2658[152], tmp2658[151], tmp2658[150], tmp2658[149], tmp2658[148], tmp2658[147], tmp2658[146], tmp2658[145], tmp2658[144], tmp2658[143], tmp2658[142], tmp2658[141], tmp2658[140], tmp2658[139], tmp2658[138], tmp2658[137], tmp2658[136], tmp2658[135], tmp2658[134], tmp2658[133], tmp2658[132], tmp2658[131], tmp2658[130], tmp2658[129], tmp2658[128], tmp2658[127], tmp2658[126], tmp2658[125], tmp2658[124], tmp2658[123], tmp2658[122], tmp2658[121], tmp2658[120], tmp2658[119], tmp2658[118], tmp2658[117], tmp2658[116], tmp2658[115], tmp2658[114], tmp2658[113], tmp2658[112], tmp2658[111], tmp2658[110], tmp2658[109], tmp2658[108], tmp2658[107], tmp2658[106], tmp2658[105], tmp2658[104], tmp2658[103], tmp2658[102], tmp2658[101], tmp2658[100], tmp2658[99], tmp2658[98], tmp2658[97], tmp2658[96], tmp2658[95], tmp2658[94], tmp2658[93], tmp2658[92], tmp2658[91], tmp2658[90], tmp2658[89], tmp2658[88], tmp2658[87], tmp2658[86], tmp2658[85], tmp2658[84], tmp2658[83], tmp2658[82], tmp2658[81], tmp2658[80], tmp2658[79], tmp2658[78], tmp2658[77], tmp2658[76], tmp2658[75], tmp2658[74], tmp2658[73], tmp2658[72], tmp2658[71], tmp2658[70], tmp2658[69], tmp2658[68], tmp2658[67], tmp2658[66], tmp2658[65], tmp2658[64], tmp2658[63], tmp2658[62], tmp2658[61], tmp2658[60], tmp2658[59], tmp2658[58], tmp2658[57], tmp2658[56], tmp2658[55], tmp2658[54], tmp2658[53], tmp2658[52], tmp2658[51], tmp2658[50], tmp2658[49], tmp2658[48], tmp2658[47], tmp2658[46], tmp2658[45], tmp2658[44], tmp2658[43], tmp2658[42], tmp2658[41], tmp2658[40], tmp2658[39], tmp2658[38], tmp2658[37], tmp2658[36], tmp2658[35], tmp2658[34], tmp2658[33], tmp2658[32], tmp2658[31], tmp2658[30], tmp2658[29], tmp2658[28], tmp2658[27], tmp2658[26], tmp2658[25], tmp2658[24], tmp2658[23], tmp2658[22], tmp2658[21], tmp2658[20], tmp2658[19], tmp2658[18], tmp2658[17], tmp2658[16], tmp2658[15], tmp2658[14], tmp2658[13], tmp2658[12], tmp2658[11], tmp2658[10], tmp2658[9], tmp2658[8], tmp2658[7], tmp2658[6], tmp2658[5], tmp2658[4], tmp2658[3], tmp2658[2], tmp2658[1], tmp2658[0]};
    assign tmp2660 = ~tmp35;
    assign tmp2661 = ~tmp36;
    assign tmp2662 = tmp2660 & tmp2661;
    assign tmp2663 = ~tmp57;
    assign tmp2664 = tmp2662 & tmp2663;
    assign tmp2665 = ~tmp1034;
    assign tmp2666 = tmp2664 & tmp2665;
    assign tmp2667 = tmp2666 & tmp2071;
    assign tmp2668 = ~tmp2583;
    assign tmp2669 = tmp2667 & tmp2668;
    assign tmp2670 = tmp2669 & tmp23;
    assign tmp2671 = tmp2670 & tmp2627;
    assign tmp2672 = tmp12 == _ver_out_tmp_65;
    assign tmp2673 = {const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0, const_304_0};
    assign tmp2674 = {tmp2673, const_303_0};
    assign tmp2675 = tmp2674 - tmp12;
    assign tmp2676 = {const_306_0, const_306_0};
    assign tmp2677 = {tmp2676, const_305_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp2678 = tmp2672 ? tmp2677 : tmp2675;
    assign tmp2679 = {tmp2678[255], tmp2678[254], tmp2678[253], tmp2678[252], tmp2678[251], tmp2678[250], tmp2678[249], tmp2678[248], tmp2678[247], tmp2678[246], tmp2678[245], tmp2678[244], tmp2678[243], tmp2678[242], tmp2678[241], tmp2678[240], tmp2678[239], tmp2678[238], tmp2678[237], tmp2678[236], tmp2678[235], tmp2678[234], tmp2678[233], tmp2678[232], tmp2678[231], tmp2678[230], tmp2678[229], tmp2678[228], tmp2678[227], tmp2678[226], tmp2678[225], tmp2678[224], tmp2678[223], tmp2678[222], tmp2678[221], tmp2678[220], tmp2678[219], tmp2678[218], tmp2678[217], tmp2678[216], tmp2678[215], tmp2678[214], tmp2678[213], tmp2678[212], tmp2678[211], tmp2678[210], tmp2678[209], tmp2678[208], tmp2678[207], tmp2678[206], tmp2678[205], tmp2678[204], tmp2678[203], tmp2678[202], tmp2678[201], tmp2678[200], tmp2678[199], tmp2678[198], tmp2678[197], tmp2678[196], tmp2678[195], tmp2678[194], tmp2678[193], tmp2678[192], tmp2678[191], tmp2678[190], tmp2678[189], tmp2678[188], tmp2678[187], tmp2678[186], tmp2678[185], tmp2678[184], tmp2678[183], tmp2678[182], tmp2678[181], tmp2678[180], tmp2678[179], tmp2678[178], tmp2678[177], tmp2678[176], tmp2678[175], tmp2678[174], tmp2678[173], tmp2678[172], tmp2678[171], tmp2678[170], tmp2678[169], tmp2678[168], tmp2678[167], tmp2678[166], tmp2678[165], tmp2678[164], tmp2678[163], tmp2678[162], tmp2678[161], tmp2678[160], tmp2678[159], tmp2678[158], tmp2678[157], tmp2678[156], tmp2678[155], tmp2678[154], tmp2678[153], tmp2678[152], tmp2678[151], tmp2678[150], tmp2678[149], tmp2678[148], tmp2678[147], tmp2678[146], tmp2678[145], tmp2678[144], tmp2678[143], tmp2678[142], tmp2678[141], tmp2678[140], tmp2678[139], tmp2678[138], tmp2678[137], tmp2678[136], tmp2678[135], tmp2678[134], tmp2678[133], tmp2678[132], tmp2678[131], tmp2678[130], tmp2678[129], tmp2678[128], tmp2678[127], tmp2678[126], tmp2678[125], tmp2678[124], tmp2678[123], tmp2678[122], tmp2678[121], tmp2678[120], tmp2678[119], tmp2678[118], tmp2678[117], tmp2678[116], tmp2678[115], tmp2678[114], tmp2678[113], tmp2678[112], tmp2678[111], tmp2678[110], tmp2678[109], tmp2678[108], tmp2678[107], tmp2678[106], tmp2678[105], tmp2678[104], tmp2678[103], tmp2678[102], tmp2678[101], tmp2678[100], tmp2678[99], tmp2678[98], tmp2678[97], tmp2678[96], tmp2678[95], tmp2678[94], tmp2678[93], tmp2678[92], tmp2678[91], tmp2678[90], tmp2678[89], tmp2678[88], tmp2678[87], tmp2678[86], tmp2678[85], tmp2678[84], tmp2678[83], tmp2678[82], tmp2678[81], tmp2678[80], tmp2678[79], tmp2678[78], tmp2678[77], tmp2678[76], tmp2678[75], tmp2678[74], tmp2678[73], tmp2678[72], tmp2678[71], tmp2678[70], tmp2678[69], tmp2678[68], tmp2678[67], tmp2678[66], tmp2678[65], tmp2678[64], tmp2678[63], tmp2678[62], tmp2678[61], tmp2678[60], tmp2678[59], tmp2678[58], tmp2678[57], tmp2678[56], tmp2678[55], tmp2678[54], tmp2678[53], tmp2678[52], tmp2678[51], tmp2678[50], tmp2678[49], tmp2678[48], tmp2678[47], tmp2678[46], tmp2678[45], tmp2678[44], tmp2678[43], tmp2678[42], tmp2678[41], tmp2678[40], tmp2678[39], tmp2678[38], tmp2678[37], tmp2678[36], tmp2678[35], tmp2678[34], tmp2678[33], tmp2678[32], tmp2678[31], tmp2678[30], tmp2678[29], tmp2678[28], tmp2678[27], tmp2678[26], tmp2678[25], tmp2678[24], tmp2678[23], tmp2678[22], tmp2678[21], tmp2678[20], tmp2678[19], tmp2678[18], tmp2678[17], tmp2678[16], tmp2678[15], tmp2678[14], tmp2678[13], tmp2678[12], tmp2678[11], tmp2678[10], tmp2678[9], tmp2678[8], tmp2678[7], tmp2678[6], tmp2678[5], tmp2678[4], tmp2678[3], tmp2678[2], tmp2678[1], tmp2678[0]};
    assign tmp2680 = ~tmp35;
    assign tmp2681 = ~tmp36;
    assign tmp2682 = tmp2680 & tmp2681;
    assign tmp2683 = ~tmp57;
    assign tmp2684 = tmp2682 & tmp2683;
    assign tmp2685 = ~tmp1034;
    assign tmp2686 = tmp2684 & tmp2685;
    assign tmp2687 = tmp2686 & tmp2071;
    assign tmp2688 = ~tmp2583;
    assign tmp2689 = tmp2687 & tmp2688;
    assign tmp2690 = tmp2689 & tmp23;
    assign tmp2691 = tmp2690 & tmp2627;
    assign tmp2692 = tmp13 == _ver_out_tmp_53;
    assign tmp2693 = {const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0, const_309_0};
    assign tmp2694 = {tmp2693, const_308_0};
    assign tmp2695 = tmp2694 - tmp13;
    assign tmp2696 = {const_311_0, const_311_0};
    assign tmp2697 = {tmp2696, const_310_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp2698 = tmp2692 ? tmp2697 : tmp2695;
    assign tmp2699 = {tmp2698[255], tmp2698[254], tmp2698[253], tmp2698[252], tmp2698[251], tmp2698[250], tmp2698[249], tmp2698[248], tmp2698[247], tmp2698[246], tmp2698[245], tmp2698[244], tmp2698[243], tmp2698[242], tmp2698[241], tmp2698[240], tmp2698[239], tmp2698[238], tmp2698[237], tmp2698[236], tmp2698[235], tmp2698[234], tmp2698[233], tmp2698[232], tmp2698[231], tmp2698[230], tmp2698[229], tmp2698[228], tmp2698[227], tmp2698[226], tmp2698[225], tmp2698[224], tmp2698[223], tmp2698[222], tmp2698[221], tmp2698[220], tmp2698[219], tmp2698[218], tmp2698[217], tmp2698[216], tmp2698[215], tmp2698[214], tmp2698[213], tmp2698[212], tmp2698[211], tmp2698[210], tmp2698[209], tmp2698[208], tmp2698[207], tmp2698[206], tmp2698[205], tmp2698[204], tmp2698[203], tmp2698[202], tmp2698[201], tmp2698[200], tmp2698[199], tmp2698[198], tmp2698[197], tmp2698[196], tmp2698[195], tmp2698[194], tmp2698[193], tmp2698[192], tmp2698[191], tmp2698[190], tmp2698[189], tmp2698[188], tmp2698[187], tmp2698[186], tmp2698[185], tmp2698[184], tmp2698[183], tmp2698[182], tmp2698[181], tmp2698[180], tmp2698[179], tmp2698[178], tmp2698[177], tmp2698[176], tmp2698[175], tmp2698[174], tmp2698[173], tmp2698[172], tmp2698[171], tmp2698[170], tmp2698[169], tmp2698[168], tmp2698[167], tmp2698[166], tmp2698[165], tmp2698[164], tmp2698[163], tmp2698[162], tmp2698[161], tmp2698[160], tmp2698[159], tmp2698[158], tmp2698[157], tmp2698[156], tmp2698[155], tmp2698[154], tmp2698[153], tmp2698[152], tmp2698[151], tmp2698[150], tmp2698[149], tmp2698[148], tmp2698[147], tmp2698[146], tmp2698[145], tmp2698[144], tmp2698[143], tmp2698[142], tmp2698[141], tmp2698[140], tmp2698[139], tmp2698[138], tmp2698[137], tmp2698[136], tmp2698[135], tmp2698[134], tmp2698[133], tmp2698[132], tmp2698[131], tmp2698[130], tmp2698[129], tmp2698[128], tmp2698[127], tmp2698[126], tmp2698[125], tmp2698[124], tmp2698[123], tmp2698[122], tmp2698[121], tmp2698[120], tmp2698[119], tmp2698[118], tmp2698[117], tmp2698[116], tmp2698[115], tmp2698[114], tmp2698[113], tmp2698[112], tmp2698[111], tmp2698[110], tmp2698[109], tmp2698[108], tmp2698[107], tmp2698[106], tmp2698[105], tmp2698[104], tmp2698[103], tmp2698[102], tmp2698[101], tmp2698[100], tmp2698[99], tmp2698[98], tmp2698[97], tmp2698[96], tmp2698[95], tmp2698[94], tmp2698[93], tmp2698[92], tmp2698[91], tmp2698[90], tmp2698[89], tmp2698[88], tmp2698[87], tmp2698[86], tmp2698[85], tmp2698[84], tmp2698[83], tmp2698[82], tmp2698[81], tmp2698[80], tmp2698[79], tmp2698[78], tmp2698[77], tmp2698[76], tmp2698[75], tmp2698[74], tmp2698[73], tmp2698[72], tmp2698[71], tmp2698[70], tmp2698[69], tmp2698[68], tmp2698[67], tmp2698[66], tmp2698[65], tmp2698[64], tmp2698[63], tmp2698[62], tmp2698[61], tmp2698[60], tmp2698[59], tmp2698[58], tmp2698[57], tmp2698[56], tmp2698[55], tmp2698[54], tmp2698[53], tmp2698[52], tmp2698[51], tmp2698[50], tmp2698[49], tmp2698[48], tmp2698[47], tmp2698[46], tmp2698[45], tmp2698[44], tmp2698[43], tmp2698[42], tmp2698[41], tmp2698[40], tmp2698[39], tmp2698[38], tmp2698[37], tmp2698[36], tmp2698[35], tmp2698[34], tmp2698[33], tmp2698[32], tmp2698[31], tmp2698[30], tmp2698[29], tmp2698[28], tmp2698[27], tmp2698[26], tmp2698[25], tmp2698[24], tmp2698[23], tmp2698[22], tmp2698[21], tmp2698[20], tmp2698[19], tmp2698[18], tmp2698[17], tmp2698[16], tmp2698[15], tmp2698[14], tmp2698[13], tmp2698[12], tmp2698[11], tmp2698[10], tmp2698[9], tmp2698[8], tmp2698[7], tmp2698[6], tmp2698[5], tmp2698[4], tmp2698[3], tmp2698[2], tmp2698[1], tmp2698[0]};
    assign tmp2700 = ~tmp35;
    assign tmp2701 = ~tmp36;
    assign tmp2702 = tmp2700 & tmp2701;
    assign tmp2703 = ~tmp57;
    assign tmp2704 = tmp2702 & tmp2703;
    assign tmp2705 = ~tmp1034;
    assign tmp2706 = tmp2704 & tmp2705;
    assign tmp2707 = tmp2706 & tmp2071;
    assign tmp2708 = ~tmp2583;
    assign tmp2709 = tmp2707 & tmp2708;
    assign tmp2710 = tmp2709 & tmp23;
    assign tmp2711 = tmp2710 & tmp2627;
    assign tmp2712 = tmp14 == _ver_out_tmp_66;
    assign tmp2713 = {const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0, const_314_0};
    assign tmp2714 = {tmp2713, const_313_0};
    assign tmp2715 = tmp2714 - tmp14;
    assign tmp2716 = {const_316_0, const_316_0};
    assign tmp2717 = {tmp2716, const_315_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp2718 = tmp2712 ? tmp2717 : tmp2715;
    assign tmp2719 = {tmp2718[255], tmp2718[254], tmp2718[253], tmp2718[252], tmp2718[251], tmp2718[250], tmp2718[249], tmp2718[248], tmp2718[247], tmp2718[246], tmp2718[245], tmp2718[244], tmp2718[243], tmp2718[242], tmp2718[241], tmp2718[240], tmp2718[239], tmp2718[238], tmp2718[237], tmp2718[236], tmp2718[235], tmp2718[234], tmp2718[233], tmp2718[232], tmp2718[231], tmp2718[230], tmp2718[229], tmp2718[228], tmp2718[227], tmp2718[226], tmp2718[225], tmp2718[224], tmp2718[223], tmp2718[222], tmp2718[221], tmp2718[220], tmp2718[219], tmp2718[218], tmp2718[217], tmp2718[216], tmp2718[215], tmp2718[214], tmp2718[213], tmp2718[212], tmp2718[211], tmp2718[210], tmp2718[209], tmp2718[208], tmp2718[207], tmp2718[206], tmp2718[205], tmp2718[204], tmp2718[203], tmp2718[202], tmp2718[201], tmp2718[200], tmp2718[199], tmp2718[198], tmp2718[197], tmp2718[196], tmp2718[195], tmp2718[194], tmp2718[193], tmp2718[192], tmp2718[191], tmp2718[190], tmp2718[189], tmp2718[188], tmp2718[187], tmp2718[186], tmp2718[185], tmp2718[184], tmp2718[183], tmp2718[182], tmp2718[181], tmp2718[180], tmp2718[179], tmp2718[178], tmp2718[177], tmp2718[176], tmp2718[175], tmp2718[174], tmp2718[173], tmp2718[172], tmp2718[171], tmp2718[170], tmp2718[169], tmp2718[168], tmp2718[167], tmp2718[166], tmp2718[165], tmp2718[164], tmp2718[163], tmp2718[162], tmp2718[161], tmp2718[160], tmp2718[159], tmp2718[158], tmp2718[157], tmp2718[156], tmp2718[155], tmp2718[154], tmp2718[153], tmp2718[152], tmp2718[151], tmp2718[150], tmp2718[149], tmp2718[148], tmp2718[147], tmp2718[146], tmp2718[145], tmp2718[144], tmp2718[143], tmp2718[142], tmp2718[141], tmp2718[140], tmp2718[139], tmp2718[138], tmp2718[137], tmp2718[136], tmp2718[135], tmp2718[134], tmp2718[133], tmp2718[132], tmp2718[131], tmp2718[130], tmp2718[129], tmp2718[128], tmp2718[127], tmp2718[126], tmp2718[125], tmp2718[124], tmp2718[123], tmp2718[122], tmp2718[121], tmp2718[120], tmp2718[119], tmp2718[118], tmp2718[117], tmp2718[116], tmp2718[115], tmp2718[114], tmp2718[113], tmp2718[112], tmp2718[111], tmp2718[110], tmp2718[109], tmp2718[108], tmp2718[107], tmp2718[106], tmp2718[105], tmp2718[104], tmp2718[103], tmp2718[102], tmp2718[101], tmp2718[100], tmp2718[99], tmp2718[98], tmp2718[97], tmp2718[96], tmp2718[95], tmp2718[94], tmp2718[93], tmp2718[92], tmp2718[91], tmp2718[90], tmp2718[89], tmp2718[88], tmp2718[87], tmp2718[86], tmp2718[85], tmp2718[84], tmp2718[83], tmp2718[82], tmp2718[81], tmp2718[80], tmp2718[79], tmp2718[78], tmp2718[77], tmp2718[76], tmp2718[75], tmp2718[74], tmp2718[73], tmp2718[72], tmp2718[71], tmp2718[70], tmp2718[69], tmp2718[68], tmp2718[67], tmp2718[66], tmp2718[65], tmp2718[64], tmp2718[63], tmp2718[62], tmp2718[61], tmp2718[60], tmp2718[59], tmp2718[58], tmp2718[57], tmp2718[56], tmp2718[55], tmp2718[54], tmp2718[53], tmp2718[52], tmp2718[51], tmp2718[50], tmp2718[49], tmp2718[48], tmp2718[47], tmp2718[46], tmp2718[45], tmp2718[44], tmp2718[43], tmp2718[42], tmp2718[41], tmp2718[40], tmp2718[39], tmp2718[38], tmp2718[37], tmp2718[36], tmp2718[35], tmp2718[34], tmp2718[33], tmp2718[32], tmp2718[31], tmp2718[30], tmp2718[29], tmp2718[28], tmp2718[27], tmp2718[26], tmp2718[25], tmp2718[24], tmp2718[23], tmp2718[22], tmp2718[21], tmp2718[20], tmp2718[19], tmp2718[18], tmp2718[17], tmp2718[16], tmp2718[15], tmp2718[14], tmp2718[13], tmp2718[12], tmp2718[11], tmp2718[10], tmp2718[9], tmp2718[8], tmp2718[7], tmp2718[6], tmp2718[5], tmp2718[4], tmp2718[3], tmp2718[2], tmp2718[1], tmp2718[0]};
    assign tmp2720 = ~tmp35;
    assign tmp2721 = ~tmp36;
    assign tmp2722 = tmp2720 & tmp2721;
    assign tmp2723 = ~tmp57;
    assign tmp2724 = tmp2722 & tmp2723;
    assign tmp2725 = ~tmp1034;
    assign tmp2726 = tmp2724 & tmp2725;
    assign tmp2727 = tmp2726 & tmp2071;
    assign tmp2728 = ~tmp2583;
    assign tmp2729 = tmp2727 & tmp2728;
    assign tmp2730 = tmp2729 & tmp23;
    assign tmp2731 = tmp2730 & tmp2627;
    assign tmp2732 = {tmp25[255], tmp25[254], tmp25[253], tmp25[252], tmp25[251], tmp25[250], tmp25[249], tmp25[248], tmp25[247], tmp25[246], tmp25[245], tmp25[244], tmp25[243], tmp25[242], tmp25[241], tmp25[240], tmp25[239], tmp25[238], tmp25[237], tmp25[236], tmp25[235], tmp25[234], tmp25[233], tmp25[232], tmp25[231], tmp25[230], tmp25[229], tmp25[228], tmp25[227], tmp25[226], tmp25[225], tmp25[224], tmp25[223], tmp25[222], tmp25[221], tmp25[220], tmp25[219], tmp25[218], tmp25[217], tmp25[216], tmp25[215], tmp25[214], tmp25[213], tmp25[212], tmp25[211], tmp25[210], tmp25[209], tmp25[208], tmp25[207], tmp25[206], tmp25[205], tmp25[204], tmp25[203], tmp25[202], tmp25[201], tmp25[200], tmp25[199], tmp25[198], tmp25[197], tmp25[196], tmp25[195], tmp25[194], tmp25[193], tmp25[192], tmp25[191], tmp25[190], tmp25[189], tmp25[188], tmp25[187], tmp25[186], tmp25[185], tmp25[184], tmp25[183], tmp25[182], tmp25[181], tmp25[180], tmp25[179], tmp25[178], tmp25[177], tmp25[176], tmp25[175], tmp25[174], tmp25[173], tmp25[172], tmp25[171], tmp25[170], tmp25[169], tmp25[168], tmp25[167], tmp25[166], tmp25[165], tmp25[164], tmp25[163], tmp25[162], tmp25[161], tmp25[160], tmp25[159], tmp25[158], tmp25[157], tmp25[156], tmp25[155], tmp25[154], tmp25[153], tmp25[152], tmp25[151], tmp25[150], tmp25[149], tmp25[148], tmp25[147], tmp25[146], tmp25[145], tmp25[144], tmp25[143], tmp25[142], tmp25[141], tmp25[140], tmp25[139], tmp25[138], tmp25[137], tmp25[136], tmp25[135], tmp25[134], tmp25[133], tmp25[132], tmp25[131], tmp25[130], tmp25[129], tmp25[128], tmp25[127], tmp25[126], tmp25[125], tmp25[124], tmp25[123], tmp25[122], tmp25[121], tmp25[120], tmp25[119], tmp25[118], tmp25[117], tmp25[116], tmp25[115], tmp25[114], tmp25[113], tmp25[112], tmp25[111], tmp25[110], tmp25[109], tmp25[108], tmp25[107], tmp25[106], tmp25[105], tmp25[104], tmp25[103], tmp25[102], tmp25[101], tmp25[100], tmp25[99], tmp25[98], tmp25[97], tmp25[96], tmp25[95], tmp25[94], tmp25[93], tmp25[92], tmp25[91], tmp25[90], tmp25[89], tmp25[88], tmp25[87], tmp25[86], tmp25[85], tmp25[84], tmp25[83], tmp25[82], tmp25[81], tmp25[80], tmp25[79], tmp25[78], tmp25[77], tmp25[76], tmp25[75], tmp25[74], tmp25[73], tmp25[72], tmp25[71], tmp25[70], tmp25[69], tmp25[68], tmp25[67], tmp25[66], tmp25[65], tmp25[64], tmp25[63], tmp25[62], tmp25[61], tmp25[60], tmp25[59], tmp25[58], tmp25[57], tmp25[56], tmp25[55], tmp25[54], tmp25[53], tmp25[52], tmp25[51], tmp25[50], tmp25[49], tmp25[48], tmp25[47], tmp25[46], tmp25[45], tmp25[44], tmp25[43], tmp25[42], tmp25[41], tmp25[40], tmp25[39], tmp25[38], tmp25[37], tmp25[36], tmp25[35], tmp25[34], tmp25[33], tmp25[32], tmp25[31], tmp25[30], tmp25[29], tmp25[28], tmp25[27], tmp25[26], tmp25[25], tmp25[24], tmp25[23], tmp25[22], tmp25[21], tmp25[20], tmp25[19], tmp25[18], tmp25[17], tmp25[16], tmp25[15], tmp25[14], tmp25[13], tmp25[12], tmp25[11], tmp25[10], tmp25[9], tmp25[8], tmp25[7], tmp25[6], tmp25[5], tmp25[4], tmp25[3], tmp25[2], tmp25[1]};
    assign tmp2733 = {tmp2732[254]};
    assign tmp2734 = {tmp2733};
    assign tmp2735 = {tmp2734, tmp2732};
    assign tmp2736 = {tmp2735[255]};
    assign tmp2737 = {tmp29[255]};
    assign tmp2738 = tmp29 - tmp2735;
    assign tmp2739 = {tmp2738[256]};
    assign tmp2740 = {tmp2735[255]};
    assign tmp2741 = ~tmp2740;
    assign tmp2742 = tmp2739 ^ tmp2741;
    assign tmp2743 = {tmp29[255]};
    assign tmp2744 = ~tmp2743;
    assign tmp2745 = tmp2742 ^ tmp2744;
    assign tmp2746 = tmp2735 == tmp29;
    assign tmp2747 = tmp2745 | tmp2746;
    assign tmp2748 = {tmp26[255], tmp26[254], tmp26[253], tmp26[252], tmp26[251], tmp26[250], tmp26[249], tmp26[248], tmp26[247], tmp26[246], tmp26[245], tmp26[244], tmp26[243], tmp26[242], tmp26[241], tmp26[240], tmp26[239], tmp26[238], tmp26[237], tmp26[236], tmp26[235], tmp26[234], tmp26[233], tmp26[232], tmp26[231], tmp26[230], tmp26[229], tmp26[228], tmp26[227], tmp26[226], tmp26[225], tmp26[224], tmp26[223], tmp26[222], tmp26[221], tmp26[220], tmp26[219], tmp26[218], tmp26[217], tmp26[216], tmp26[215], tmp26[214], tmp26[213], tmp26[212], tmp26[211], tmp26[210], tmp26[209], tmp26[208], tmp26[207], tmp26[206], tmp26[205], tmp26[204], tmp26[203], tmp26[202], tmp26[201], tmp26[200], tmp26[199], tmp26[198], tmp26[197], tmp26[196], tmp26[195], tmp26[194], tmp26[193], tmp26[192], tmp26[191], tmp26[190], tmp26[189], tmp26[188], tmp26[187], tmp26[186], tmp26[185], tmp26[184], tmp26[183], tmp26[182], tmp26[181], tmp26[180], tmp26[179], tmp26[178], tmp26[177], tmp26[176], tmp26[175], tmp26[174], tmp26[173], tmp26[172], tmp26[171], tmp26[170], tmp26[169], tmp26[168], tmp26[167], tmp26[166], tmp26[165], tmp26[164], tmp26[163], tmp26[162], tmp26[161], tmp26[160], tmp26[159], tmp26[158], tmp26[157], tmp26[156], tmp26[155], tmp26[154], tmp26[153], tmp26[152], tmp26[151], tmp26[150], tmp26[149], tmp26[148], tmp26[147], tmp26[146], tmp26[145], tmp26[144], tmp26[143], tmp26[142], tmp26[141], tmp26[140], tmp26[139], tmp26[138], tmp26[137], tmp26[136], tmp26[135], tmp26[134], tmp26[133], tmp26[132], tmp26[131], tmp26[130], tmp26[129], tmp26[128], tmp26[127], tmp26[126], tmp26[125], tmp26[124], tmp26[123], tmp26[122], tmp26[121], tmp26[120], tmp26[119], tmp26[118], tmp26[117], tmp26[116], tmp26[115], tmp26[114], tmp26[113], tmp26[112], tmp26[111], tmp26[110], tmp26[109], tmp26[108], tmp26[107], tmp26[106], tmp26[105], tmp26[104], tmp26[103], tmp26[102], tmp26[101], tmp26[100], tmp26[99], tmp26[98], tmp26[97], tmp26[96], tmp26[95], tmp26[94], tmp26[93], tmp26[92], tmp26[91], tmp26[90], tmp26[89], tmp26[88], tmp26[87], tmp26[86], tmp26[85], tmp26[84], tmp26[83], tmp26[82], tmp26[81], tmp26[80], tmp26[79], tmp26[78], tmp26[77], tmp26[76], tmp26[75], tmp26[74], tmp26[73], tmp26[72], tmp26[71], tmp26[70], tmp26[69], tmp26[68], tmp26[67], tmp26[66], tmp26[65], tmp26[64], tmp26[63], tmp26[62], tmp26[61], tmp26[60], tmp26[59], tmp26[58], tmp26[57], tmp26[56], tmp26[55], tmp26[54], tmp26[53], tmp26[52], tmp26[51], tmp26[50], tmp26[49], tmp26[48], tmp26[47], tmp26[46], tmp26[45], tmp26[44], tmp26[43], tmp26[42], tmp26[41], tmp26[40], tmp26[39], tmp26[38], tmp26[37], tmp26[36], tmp26[35], tmp26[34], tmp26[33], tmp26[32], tmp26[31], tmp26[30], tmp26[29], tmp26[28], tmp26[27], tmp26[26], tmp26[25], tmp26[24], tmp26[23], tmp26[22], tmp26[21], tmp26[20], tmp26[19], tmp26[18], tmp26[17], tmp26[16], tmp26[15], tmp26[14], tmp26[13], tmp26[12], tmp26[11], tmp26[10], tmp26[9], tmp26[8], tmp26[7], tmp26[6], tmp26[5], tmp26[4], tmp26[3], tmp26[2], tmp26[1]};
    assign tmp2749 = {tmp2748[254]};
    assign tmp2750 = {tmp2749};
    assign tmp2751 = {tmp2750, tmp2748};
    assign tmp2752 = {tmp2751[255]};
    assign tmp2753 = {tmp30[255]};
    assign tmp2754 = tmp30 - tmp2751;
    assign tmp2755 = {tmp2754[256]};
    assign tmp2756 = {tmp2751[255]};
    assign tmp2757 = ~tmp2756;
    assign tmp2758 = tmp2755 ^ tmp2757;
    assign tmp2759 = {tmp30[255]};
    assign tmp2760 = ~tmp2759;
    assign tmp2761 = tmp2758 ^ tmp2760;
    assign tmp2762 = tmp2751 == tmp30;
    assign tmp2763 = tmp2761 | tmp2762;
    assign tmp2764 = tmp2747 & tmp2763;
    assign tmp2765 = {tmp27[255], tmp27[254], tmp27[253], tmp27[252], tmp27[251], tmp27[250], tmp27[249], tmp27[248], tmp27[247], tmp27[246], tmp27[245], tmp27[244], tmp27[243], tmp27[242], tmp27[241], tmp27[240], tmp27[239], tmp27[238], tmp27[237], tmp27[236], tmp27[235], tmp27[234], tmp27[233], tmp27[232], tmp27[231], tmp27[230], tmp27[229], tmp27[228], tmp27[227], tmp27[226], tmp27[225], tmp27[224], tmp27[223], tmp27[222], tmp27[221], tmp27[220], tmp27[219], tmp27[218], tmp27[217], tmp27[216], tmp27[215], tmp27[214], tmp27[213], tmp27[212], tmp27[211], tmp27[210], tmp27[209], tmp27[208], tmp27[207], tmp27[206], tmp27[205], tmp27[204], tmp27[203], tmp27[202], tmp27[201], tmp27[200], tmp27[199], tmp27[198], tmp27[197], tmp27[196], tmp27[195], tmp27[194], tmp27[193], tmp27[192], tmp27[191], tmp27[190], tmp27[189], tmp27[188], tmp27[187], tmp27[186], tmp27[185], tmp27[184], tmp27[183], tmp27[182], tmp27[181], tmp27[180], tmp27[179], tmp27[178], tmp27[177], tmp27[176], tmp27[175], tmp27[174], tmp27[173], tmp27[172], tmp27[171], tmp27[170], tmp27[169], tmp27[168], tmp27[167], tmp27[166], tmp27[165], tmp27[164], tmp27[163], tmp27[162], tmp27[161], tmp27[160], tmp27[159], tmp27[158], tmp27[157], tmp27[156], tmp27[155], tmp27[154], tmp27[153], tmp27[152], tmp27[151], tmp27[150], tmp27[149], tmp27[148], tmp27[147], tmp27[146], tmp27[145], tmp27[144], tmp27[143], tmp27[142], tmp27[141], tmp27[140], tmp27[139], tmp27[138], tmp27[137], tmp27[136], tmp27[135], tmp27[134], tmp27[133], tmp27[132], tmp27[131], tmp27[130], tmp27[129], tmp27[128], tmp27[127], tmp27[126], tmp27[125], tmp27[124], tmp27[123], tmp27[122], tmp27[121], tmp27[120], tmp27[119], tmp27[118], tmp27[117], tmp27[116], tmp27[115], tmp27[114], tmp27[113], tmp27[112], tmp27[111], tmp27[110], tmp27[109], tmp27[108], tmp27[107], tmp27[106], tmp27[105], tmp27[104], tmp27[103], tmp27[102], tmp27[101], tmp27[100], tmp27[99], tmp27[98], tmp27[97], tmp27[96], tmp27[95], tmp27[94], tmp27[93], tmp27[92], tmp27[91], tmp27[90], tmp27[89], tmp27[88], tmp27[87], tmp27[86], tmp27[85], tmp27[84], tmp27[83], tmp27[82], tmp27[81], tmp27[80], tmp27[79], tmp27[78], tmp27[77], tmp27[76], tmp27[75], tmp27[74], tmp27[73], tmp27[72], tmp27[71], tmp27[70], tmp27[69], tmp27[68], tmp27[67], tmp27[66], tmp27[65], tmp27[64], tmp27[63], tmp27[62], tmp27[61], tmp27[60], tmp27[59], tmp27[58], tmp27[57], tmp27[56], tmp27[55], tmp27[54], tmp27[53], tmp27[52], tmp27[51], tmp27[50], tmp27[49], tmp27[48], tmp27[47], tmp27[46], tmp27[45], tmp27[44], tmp27[43], tmp27[42], tmp27[41], tmp27[40], tmp27[39], tmp27[38], tmp27[37], tmp27[36], tmp27[35], tmp27[34], tmp27[33], tmp27[32], tmp27[31], tmp27[30], tmp27[29], tmp27[28], tmp27[27], tmp27[26], tmp27[25], tmp27[24], tmp27[23], tmp27[22], tmp27[21], tmp27[20], tmp27[19], tmp27[18], tmp27[17], tmp27[16], tmp27[15], tmp27[14], tmp27[13], tmp27[12], tmp27[11], tmp27[10], tmp27[9], tmp27[8], tmp27[7], tmp27[6], tmp27[5], tmp27[4], tmp27[3], tmp27[2], tmp27[1]};
    assign tmp2766 = {tmp2765[254]};
    assign tmp2767 = {tmp2766};
    assign tmp2768 = {tmp2767, tmp2765};
    assign tmp2769 = {tmp2768[255]};
    assign tmp2770 = {tmp31[255]};
    assign tmp2771 = tmp31 - tmp2768;
    assign tmp2772 = {tmp2771[256]};
    assign tmp2773 = {tmp2768[255]};
    assign tmp2774 = ~tmp2773;
    assign tmp2775 = tmp2772 ^ tmp2774;
    assign tmp2776 = {tmp31[255]};
    assign tmp2777 = ~tmp2776;
    assign tmp2778 = tmp2775 ^ tmp2777;
    assign tmp2779 = tmp2768 == tmp31;
    assign tmp2780 = tmp2778 | tmp2779;
    assign tmp2781 = tmp2764 & tmp2780;
    assign tmp2782 = {tmp28[255], tmp28[254], tmp28[253], tmp28[252], tmp28[251], tmp28[250], tmp28[249], tmp28[248], tmp28[247], tmp28[246], tmp28[245], tmp28[244], tmp28[243], tmp28[242], tmp28[241], tmp28[240], tmp28[239], tmp28[238], tmp28[237], tmp28[236], tmp28[235], tmp28[234], tmp28[233], tmp28[232], tmp28[231], tmp28[230], tmp28[229], tmp28[228], tmp28[227], tmp28[226], tmp28[225], tmp28[224], tmp28[223], tmp28[222], tmp28[221], tmp28[220], tmp28[219], tmp28[218], tmp28[217], tmp28[216], tmp28[215], tmp28[214], tmp28[213], tmp28[212], tmp28[211], tmp28[210], tmp28[209], tmp28[208], tmp28[207], tmp28[206], tmp28[205], tmp28[204], tmp28[203], tmp28[202], tmp28[201], tmp28[200], tmp28[199], tmp28[198], tmp28[197], tmp28[196], tmp28[195], tmp28[194], tmp28[193], tmp28[192], tmp28[191], tmp28[190], tmp28[189], tmp28[188], tmp28[187], tmp28[186], tmp28[185], tmp28[184], tmp28[183], tmp28[182], tmp28[181], tmp28[180], tmp28[179], tmp28[178], tmp28[177], tmp28[176], tmp28[175], tmp28[174], tmp28[173], tmp28[172], tmp28[171], tmp28[170], tmp28[169], tmp28[168], tmp28[167], tmp28[166], tmp28[165], tmp28[164], tmp28[163], tmp28[162], tmp28[161], tmp28[160], tmp28[159], tmp28[158], tmp28[157], tmp28[156], tmp28[155], tmp28[154], tmp28[153], tmp28[152], tmp28[151], tmp28[150], tmp28[149], tmp28[148], tmp28[147], tmp28[146], tmp28[145], tmp28[144], tmp28[143], tmp28[142], tmp28[141], tmp28[140], tmp28[139], tmp28[138], tmp28[137], tmp28[136], tmp28[135], tmp28[134], tmp28[133], tmp28[132], tmp28[131], tmp28[130], tmp28[129], tmp28[128], tmp28[127], tmp28[126], tmp28[125], tmp28[124], tmp28[123], tmp28[122], tmp28[121], tmp28[120], tmp28[119], tmp28[118], tmp28[117], tmp28[116], tmp28[115], tmp28[114], tmp28[113], tmp28[112], tmp28[111], tmp28[110], tmp28[109], tmp28[108], tmp28[107], tmp28[106], tmp28[105], tmp28[104], tmp28[103], tmp28[102], tmp28[101], tmp28[100], tmp28[99], tmp28[98], tmp28[97], tmp28[96], tmp28[95], tmp28[94], tmp28[93], tmp28[92], tmp28[91], tmp28[90], tmp28[89], tmp28[88], tmp28[87], tmp28[86], tmp28[85], tmp28[84], tmp28[83], tmp28[82], tmp28[81], tmp28[80], tmp28[79], tmp28[78], tmp28[77], tmp28[76], tmp28[75], tmp28[74], tmp28[73], tmp28[72], tmp28[71], tmp28[70], tmp28[69], tmp28[68], tmp28[67], tmp28[66], tmp28[65], tmp28[64], tmp28[63], tmp28[62], tmp28[61], tmp28[60], tmp28[59], tmp28[58], tmp28[57], tmp28[56], tmp28[55], tmp28[54], tmp28[53], tmp28[52], tmp28[51], tmp28[50], tmp28[49], tmp28[48], tmp28[47], tmp28[46], tmp28[45], tmp28[44], tmp28[43], tmp28[42], tmp28[41], tmp28[40], tmp28[39], tmp28[38], tmp28[37], tmp28[36], tmp28[35], tmp28[34], tmp28[33], tmp28[32], tmp28[31], tmp28[30], tmp28[29], tmp28[28], tmp28[27], tmp28[26], tmp28[25], tmp28[24], tmp28[23], tmp28[22], tmp28[21], tmp28[20], tmp28[19], tmp28[18], tmp28[17], tmp28[16], tmp28[15], tmp28[14], tmp28[13], tmp28[12], tmp28[11], tmp28[10], tmp28[9], tmp28[8], tmp28[7], tmp28[6], tmp28[5], tmp28[4], tmp28[3], tmp28[2], tmp28[1]};
    assign tmp2783 = {tmp2782[254]};
    assign tmp2784 = {tmp2783};
    assign tmp2785 = {tmp2784, tmp2782};
    assign tmp2786 = {tmp2785[255]};
    assign tmp2787 = {tmp32[255]};
    assign tmp2788 = tmp32 - tmp2785;
    assign tmp2789 = {tmp2788[256]};
    assign tmp2790 = {tmp2785[255]};
    assign tmp2791 = ~tmp2790;
    assign tmp2792 = tmp2789 ^ tmp2791;
    assign tmp2793 = {tmp32[255]};
    assign tmp2794 = ~tmp2793;
    assign tmp2795 = tmp2792 ^ tmp2794;
    assign tmp2796 = tmp2785 == tmp32;
    assign tmp2797 = tmp2795 | tmp2796;
    assign tmp2798 = tmp2781 & tmp2797;
    assign tmp2799 = ~tmp35;
    assign tmp2800 = ~tmp36;
    assign tmp2801 = tmp2799 & tmp2800;
    assign tmp2802 = ~tmp57;
    assign tmp2803 = tmp2801 & tmp2802;
    assign tmp2804 = ~tmp1034;
    assign tmp2805 = tmp2803 & tmp2804;
    assign tmp2806 = tmp2805 & tmp2071;
    assign tmp2807 = ~tmp2583;
    assign tmp2808 = tmp2806 & tmp2807;
    assign tmp2809 = tmp2808 & tmp23;
    assign tmp2810 = ~tmp2627;
    assign tmp2811 = tmp2809 & tmp2810;
    assign tmp2812 = tmp2811 & tmp2798;
    assign tmp2813 = ~tmp35;
    assign tmp2814 = ~tmp36;
    assign tmp2815 = tmp2813 & tmp2814;
    assign tmp2816 = ~tmp57;
    assign tmp2817 = tmp2815 & tmp2816;
    assign tmp2818 = ~tmp1034;
    assign tmp2819 = tmp2817 & tmp2818;
    assign tmp2820 = tmp2819 & tmp2071;
    assign tmp2821 = ~tmp2583;
    assign tmp2822 = tmp2820 & tmp2821;
    assign tmp2823 = tmp2822 & tmp23;
    assign tmp2824 = ~tmp2627;
    assign tmp2825 = tmp2823 & tmp2824;
    assign tmp2826 = tmp2825 & tmp2798;
    assign tmp2827 = {tmp25[255], tmp25[254], tmp25[253], tmp25[252], tmp25[251], tmp25[250], tmp25[249], tmp25[248], tmp25[247], tmp25[246], tmp25[245], tmp25[244], tmp25[243], tmp25[242], tmp25[241], tmp25[240], tmp25[239], tmp25[238], tmp25[237], tmp25[236], tmp25[235], tmp25[234], tmp25[233], tmp25[232], tmp25[231], tmp25[230], tmp25[229], tmp25[228], tmp25[227], tmp25[226], tmp25[225], tmp25[224], tmp25[223], tmp25[222], tmp25[221], tmp25[220], tmp25[219], tmp25[218], tmp25[217], tmp25[216], tmp25[215], tmp25[214], tmp25[213], tmp25[212], tmp25[211], tmp25[210], tmp25[209], tmp25[208], tmp25[207], tmp25[206], tmp25[205], tmp25[204], tmp25[203], tmp25[202], tmp25[201], tmp25[200], tmp25[199], tmp25[198], tmp25[197], tmp25[196], tmp25[195], tmp25[194], tmp25[193], tmp25[192], tmp25[191], tmp25[190], tmp25[189], tmp25[188], tmp25[187], tmp25[186], tmp25[185], tmp25[184], tmp25[183], tmp25[182], tmp25[181], tmp25[180], tmp25[179], tmp25[178], tmp25[177], tmp25[176], tmp25[175], tmp25[174], tmp25[173], tmp25[172], tmp25[171], tmp25[170], tmp25[169], tmp25[168], tmp25[167], tmp25[166], tmp25[165], tmp25[164], tmp25[163], tmp25[162], tmp25[161], tmp25[160], tmp25[159], tmp25[158], tmp25[157], tmp25[156], tmp25[155], tmp25[154], tmp25[153], tmp25[152], tmp25[151], tmp25[150], tmp25[149], tmp25[148], tmp25[147], tmp25[146], tmp25[145], tmp25[144], tmp25[143], tmp25[142], tmp25[141], tmp25[140], tmp25[139], tmp25[138], tmp25[137], tmp25[136], tmp25[135], tmp25[134], tmp25[133], tmp25[132], tmp25[131], tmp25[130], tmp25[129], tmp25[128], tmp25[127], tmp25[126], tmp25[125], tmp25[124], tmp25[123], tmp25[122], tmp25[121], tmp25[120], tmp25[119], tmp25[118], tmp25[117], tmp25[116], tmp25[115], tmp25[114], tmp25[113], tmp25[112], tmp25[111], tmp25[110], tmp25[109], tmp25[108], tmp25[107], tmp25[106], tmp25[105], tmp25[104], tmp25[103], tmp25[102], tmp25[101], tmp25[100], tmp25[99], tmp25[98], tmp25[97], tmp25[96], tmp25[95], tmp25[94], tmp25[93], tmp25[92], tmp25[91], tmp25[90], tmp25[89], tmp25[88], tmp25[87], tmp25[86], tmp25[85], tmp25[84], tmp25[83], tmp25[82], tmp25[81], tmp25[80], tmp25[79], tmp25[78], tmp25[77], tmp25[76], tmp25[75], tmp25[74], tmp25[73], tmp25[72], tmp25[71], tmp25[70], tmp25[69], tmp25[68], tmp25[67], tmp25[66], tmp25[65], tmp25[64], tmp25[63], tmp25[62], tmp25[61], tmp25[60], tmp25[59], tmp25[58], tmp25[57], tmp25[56], tmp25[55], tmp25[54], tmp25[53], tmp25[52], tmp25[51], tmp25[50], tmp25[49], tmp25[48], tmp25[47], tmp25[46], tmp25[45], tmp25[44], tmp25[43], tmp25[42], tmp25[41], tmp25[40], tmp25[39], tmp25[38], tmp25[37], tmp25[36], tmp25[35], tmp25[34], tmp25[33], tmp25[32], tmp25[31], tmp25[30], tmp25[29], tmp25[28], tmp25[27], tmp25[26], tmp25[25], tmp25[24], tmp25[23], tmp25[22], tmp25[21], tmp25[20], tmp25[19], tmp25[18], tmp25[17], tmp25[16], tmp25[15], tmp25[14], tmp25[13], tmp25[12], tmp25[11], tmp25[10], tmp25[9], tmp25[8], tmp25[7], tmp25[6], tmp25[5], tmp25[4], tmp25[3], tmp25[2], tmp25[1]};
    assign tmp2828 = {tmp2827[254]};
    assign tmp2829 = {tmp2828};
    assign tmp2830 = {tmp2829, tmp2827};
    assign tmp2831 = ~tmp35;
    assign tmp2832 = ~tmp36;
    assign tmp2833 = tmp2831 & tmp2832;
    assign tmp2834 = ~tmp57;
    assign tmp2835 = tmp2833 & tmp2834;
    assign tmp2836 = ~tmp1034;
    assign tmp2837 = tmp2835 & tmp2836;
    assign tmp2838 = tmp2837 & tmp2071;
    assign tmp2839 = ~tmp2583;
    assign tmp2840 = tmp2838 & tmp2839;
    assign tmp2841 = tmp2840 & tmp23;
    assign tmp2842 = ~tmp2627;
    assign tmp2843 = tmp2841 & tmp2842;
    assign tmp2844 = tmp2843 & tmp2798;
    assign tmp2845 = tmp2844 & tmp24;
    assign tmp2846 = {tmp26[255], tmp26[254], tmp26[253], tmp26[252], tmp26[251], tmp26[250], tmp26[249], tmp26[248], tmp26[247], tmp26[246], tmp26[245], tmp26[244], tmp26[243], tmp26[242], tmp26[241], tmp26[240], tmp26[239], tmp26[238], tmp26[237], tmp26[236], tmp26[235], tmp26[234], tmp26[233], tmp26[232], tmp26[231], tmp26[230], tmp26[229], tmp26[228], tmp26[227], tmp26[226], tmp26[225], tmp26[224], tmp26[223], tmp26[222], tmp26[221], tmp26[220], tmp26[219], tmp26[218], tmp26[217], tmp26[216], tmp26[215], tmp26[214], tmp26[213], tmp26[212], tmp26[211], tmp26[210], tmp26[209], tmp26[208], tmp26[207], tmp26[206], tmp26[205], tmp26[204], tmp26[203], tmp26[202], tmp26[201], tmp26[200], tmp26[199], tmp26[198], tmp26[197], tmp26[196], tmp26[195], tmp26[194], tmp26[193], tmp26[192], tmp26[191], tmp26[190], tmp26[189], tmp26[188], tmp26[187], tmp26[186], tmp26[185], tmp26[184], tmp26[183], tmp26[182], tmp26[181], tmp26[180], tmp26[179], tmp26[178], tmp26[177], tmp26[176], tmp26[175], tmp26[174], tmp26[173], tmp26[172], tmp26[171], tmp26[170], tmp26[169], tmp26[168], tmp26[167], tmp26[166], tmp26[165], tmp26[164], tmp26[163], tmp26[162], tmp26[161], tmp26[160], tmp26[159], tmp26[158], tmp26[157], tmp26[156], tmp26[155], tmp26[154], tmp26[153], tmp26[152], tmp26[151], tmp26[150], tmp26[149], tmp26[148], tmp26[147], tmp26[146], tmp26[145], tmp26[144], tmp26[143], tmp26[142], tmp26[141], tmp26[140], tmp26[139], tmp26[138], tmp26[137], tmp26[136], tmp26[135], tmp26[134], tmp26[133], tmp26[132], tmp26[131], tmp26[130], tmp26[129], tmp26[128], tmp26[127], tmp26[126], tmp26[125], tmp26[124], tmp26[123], tmp26[122], tmp26[121], tmp26[120], tmp26[119], tmp26[118], tmp26[117], tmp26[116], tmp26[115], tmp26[114], tmp26[113], tmp26[112], tmp26[111], tmp26[110], tmp26[109], tmp26[108], tmp26[107], tmp26[106], tmp26[105], tmp26[104], tmp26[103], tmp26[102], tmp26[101], tmp26[100], tmp26[99], tmp26[98], tmp26[97], tmp26[96], tmp26[95], tmp26[94], tmp26[93], tmp26[92], tmp26[91], tmp26[90], tmp26[89], tmp26[88], tmp26[87], tmp26[86], tmp26[85], tmp26[84], tmp26[83], tmp26[82], tmp26[81], tmp26[80], tmp26[79], tmp26[78], tmp26[77], tmp26[76], tmp26[75], tmp26[74], tmp26[73], tmp26[72], tmp26[71], tmp26[70], tmp26[69], tmp26[68], tmp26[67], tmp26[66], tmp26[65], tmp26[64], tmp26[63], tmp26[62], tmp26[61], tmp26[60], tmp26[59], tmp26[58], tmp26[57], tmp26[56], tmp26[55], tmp26[54], tmp26[53], tmp26[52], tmp26[51], tmp26[50], tmp26[49], tmp26[48], tmp26[47], tmp26[46], tmp26[45], tmp26[44], tmp26[43], tmp26[42], tmp26[41], tmp26[40], tmp26[39], tmp26[38], tmp26[37], tmp26[36], tmp26[35], tmp26[34], tmp26[33], tmp26[32], tmp26[31], tmp26[30], tmp26[29], tmp26[28], tmp26[27], tmp26[26], tmp26[25], tmp26[24], tmp26[23], tmp26[22], tmp26[21], tmp26[20], tmp26[19], tmp26[18], tmp26[17], tmp26[16], tmp26[15], tmp26[14], tmp26[13], tmp26[12], tmp26[11], tmp26[10], tmp26[9], tmp26[8], tmp26[7], tmp26[6], tmp26[5], tmp26[4], tmp26[3], tmp26[2], tmp26[1]};
    assign tmp2847 = {tmp2846[254]};
    assign tmp2848 = {tmp2847};
    assign tmp2849 = {tmp2848, tmp2846};
    assign tmp2850 = ~tmp35;
    assign tmp2851 = ~tmp36;
    assign tmp2852 = tmp2850 & tmp2851;
    assign tmp2853 = ~tmp57;
    assign tmp2854 = tmp2852 & tmp2853;
    assign tmp2855 = ~tmp1034;
    assign tmp2856 = tmp2854 & tmp2855;
    assign tmp2857 = tmp2856 & tmp2071;
    assign tmp2858 = ~tmp2583;
    assign tmp2859 = tmp2857 & tmp2858;
    assign tmp2860 = tmp2859 & tmp23;
    assign tmp2861 = ~tmp2627;
    assign tmp2862 = tmp2860 & tmp2861;
    assign tmp2863 = tmp2862 & tmp2798;
    assign tmp2864 = tmp2863 & tmp24;
    assign tmp2865 = {tmp27[255], tmp27[254], tmp27[253], tmp27[252], tmp27[251], tmp27[250], tmp27[249], tmp27[248], tmp27[247], tmp27[246], tmp27[245], tmp27[244], tmp27[243], tmp27[242], tmp27[241], tmp27[240], tmp27[239], tmp27[238], tmp27[237], tmp27[236], tmp27[235], tmp27[234], tmp27[233], tmp27[232], tmp27[231], tmp27[230], tmp27[229], tmp27[228], tmp27[227], tmp27[226], tmp27[225], tmp27[224], tmp27[223], tmp27[222], tmp27[221], tmp27[220], tmp27[219], tmp27[218], tmp27[217], tmp27[216], tmp27[215], tmp27[214], tmp27[213], tmp27[212], tmp27[211], tmp27[210], tmp27[209], tmp27[208], tmp27[207], tmp27[206], tmp27[205], tmp27[204], tmp27[203], tmp27[202], tmp27[201], tmp27[200], tmp27[199], tmp27[198], tmp27[197], tmp27[196], tmp27[195], tmp27[194], tmp27[193], tmp27[192], tmp27[191], tmp27[190], tmp27[189], tmp27[188], tmp27[187], tmp27[186], tmp27[185], tmp27[184], tmp27[183], tmp27[182], tmp27[181], tmp27[180], tmp27[179], tmp27[178], tmp27[177], tmp27[176], tmp27[175], tmp27[174], tmp27[173], tmp27[172], tmp27[171], tmp27[170], tmp27[169], tmp27[168], tmp27[167], tmp27[166], tmp27[165], tmp27[164], tmp27[163], tmp27[162], tmp27[161], tmp27[160], tmp27[159], tmp27[158], tmp27[157], tmp27[156], tmp27[155], tmp27[154], tmp27[153], tmp27[152], tmp27[151], tmp27[150], tmp27[149], tmp27[148], tmp27[147], tmp27[146], tmp27[145], tmp27[144], tmp27[143], tmp27[142], tmp27[141], tmp27[140], tmp27[139], tmp27[138], tmp27[137], tmp27[136], tmp27[135], tmp27[134], tmp27[133], tmp27[132], tmp27[131], tmp27[130], tmp27[129], tmp27[128], tmp27[127], tmp27[126], tmp27[125], tmp27[124], tmp27[123], tmp27[122], tmp27[121], tmp27[120], tmp27[119], tmp27[118], tmp27[117], tmp27[116], tmp27[115], tmp27[114], tmp27[113], tmp27[112], tmp27[111], tmp27[110], tmp27[109], tmp27[108], tmp27[107], tmp27[106], tmp27[105], tmp27[104], tmp27[103], tmp27[102], tmp27[101], tmp27[100], tmp27[99], tmp27[98], tmp27[97], tmp27[96], tmp27[95], tmp27[94], tmp27[93], tmp27[92], tmp27[91], tmp27[90], tmp27[89], tmp27[88], tmp27[87], tmp27[86], tmp27[85], tmp27[84], tmp27[83], tmp27[82], tmp27[81], tmp27[80], tmp27[79], tmp27[78], tmp27[77], tmp27[76], tmp27[75], tmp27[74], tmp27[73], tmp27[72], tmp27[71], tmp27[70], tmp27[69], tmp27[68], tmp27[67], tmp27[66], tmp27[65], tmp27[64], tmp27[63], tmp27[62], tmp27[61], tmp27[60], tmp27[59], tmp27[58], tmp27[57], tmp27[56], tmp27[55], tmp27[54], tmp27[53], tmp27[52], tmp27[51], tmp27[50], tmp27[49], tmp27[48], tmp27[47], tmp27[46], tmp27[45], tmp27[44], tmp27[43], tmp27[42], tmp27[41], tmp27[40], tmp27[39], tmp27[38], tmp27[37], tmp27[36], tmp27[35], tmp27[34], tmp27[33], tmp27[32], tmp27[31], tmp27[30], tmp27[29], tmp27[28], tmp27[27], tmp27[26], tmp27[25], tmp27[24], tmp27[23], tmp27[22], tmp27[21], tmp27[20], tmp27[19], tmp27[18], tmp27[17], tmp27[16], tmp27[15], tmp27[14], tmp27[13], tmp27[12], tmp27[11], tmp27[10], tmp27[9], tmp27[8], tmp27[7], tmp27[6], tmp27[5], tmp27[4], tmp27[3], tmp27[2], tmp27[1]};
    assign tmp2866 = {tmp2865[254]};
    assign tmp2867 = {tmp2866};
    assign tmp2868 = {tmp2867, tmp2865};
    assign tmp2869 = ~tmp35;
    assign tmp2870 = ~tmp36;
    assign tmp2871 = tmp2869 & tmp2870;
    assign tmp2872 = ~tmp57;
    assign tmp2873 = tmp2871 & tmp2872;
    assign tmp2874 = ~tmp1034;
    assign tmp2875 = tmp2873 & tmp2874;
    assign tmp2876 = tmp2875 & tmp2071;
    assign tmp2877 = ~tmp2583;
    assign tmp2878 = tmp2876 & tmp2877;
    assign tmp2879 = tmp2878 & tmp23;
    assign tmp2880 = ~tmp2627;
    assign tmp2881 = tmp2879 & tmp2880;
    assign tmp2882 = tmp2881 & tmp2798;
    assign tmp2883 = tmp2882 & tmp24;
    assign tmp2884 = {tmp28[255], tmp28[254], tmp28[253], tmp28[252], tmp28[251], tmp28[250], tmp28[249], tmp28[248], tmp28[247], tmp28[246], tmp28[245], tmp28[244], tmp28[243], tmp28[242], tmp28[241], tmp28[240], tmp28[239], tmp28[238], tmp28[237], tmp28[236], tmp28[235], tmp28[234], tmp28[233], tmp28[232], tmp28[231], tmp28[230], tmp28[229], tmp28[228], tmp28[227], tmp28[226], tmp28[225], tmp28[224], tmp28[223], tmp28[222], tmp28[221], tmp28[220], tmp28[219], tmp28[218], tmp28[217], tmp28[216], tmp28[215], tmp28[214], tmp28[213], tmp28[212], tmp28[211], tmp28[210], tmp28[209], tmp28[208], tmp28[207], tmp28[206], tmp28[205], tmp28[204], tmp28[203], tmp28[202], tmp28[201], tmp28[200], tmp28[199], tmp28[198], tmp28[197], tmp28[196], tmp28[195], tmp28[194], tmp28[193], tmp28[192], tmp28[191], tmp28[190], tmp28[189], tmp28[188], tmp28[187], tmp28[186], tmp28[185], tmp28[184], tmp28[183], tmp28[182], tmp28[181], tmp28[180], tmp28[179], tmp28[178], tmp28[177], tmp28[176], tmp28[175], tmp28[174], tmp28[173], tmp28[172], tmp28[171], tmp28[170], tmp28[169], tmp28[168], tmp28[167], tmp28[166], tmp28[165], tmp28[164], tmp28[163], tmp28[162], tmp28[161], tmp28[160], tmp28[159], tmp28[158], tmp28[157], tmp28[156], tmp28[155], tmp28[154], tmp28[153], tmp28[152], tmp28[151], tmp28[150], tmp28[149], tmp28[148], tmp28[147], tmp28[146], tmp28[145], tmp28[144], tmp28[143], tmp28[142], tmp28[141], tmp28[140], tmp28[139], tmp28[138], tmp28[137], tmp28[136], tmp28[135], tmp28[134], tmp28[133], tmp28[132], tmp28[131], tmp28[130], tmp28[129], tmp28[128], tmp28[127], tmp28[126], tmp28[125], tmp28[124], tmp28[123], tmp28[122], tmp28[121], tmp28[120], tmp28[119], tmp28[118], tmp28[117], tmp28[116], tmp28[115], tmp28[114], tmp28[113], tmp28[112], tmp28[111], tmp28[110], tmp28[109], tmp28[108], tmp28[107], tmp28[106], tmp28[105], tmp28[104], tmp28[103], tmp28[102], tmp28[101], tmp28[100], tmp28[99], tmp28[98], tmp28[97], tmp28[96], tmp28[95], tmp28[94], tmp28[93], tmp28[92], tmp28[91], tmp28[90], tmp28[89], tmp28[88], tmp28[87], tmp28[86], tmp28[85], tmp28[84], tmp28[83], tmp28[82], tmp28[81], tmp28[80], tmp28[79], tmp28[78], tmp28[77], tmp28[76], tmp28[75], tmp28[74], tmp28[73], tmp28[72], tmp28[71], tmp28[70], tmp28[69], tmp28[68], tmp28[67], tmp28[66], tmp28[65], tmp28[64], tmp28[63], tmp28[62], tmp28[61], tmp28[60], tmp28[59], tmp28[58], tmp28[57], tmp28[56], tmp28[55], tmp28[54], tmp28[53], tmp28[52], tmp28[51], tmp28[50], tmp28[49], tmp28[48], tmp28[47], tmp28[46], tmp28[45], tmp28[44], tmp28[43], tmp28[42], tmp28[41], tmp28[40], tmp28[39], tmp28[38], tmp28[37], tmp28[36], tmp28[35], tmp28[34], tmp28[33], tmp28[32], tmp28[31], tmp28[30], tmp28[29], tmp28[28], tmp28[27], tmp28[26], tmp28[25], tmp28[24], tmp28[23], tmp28[22], tmp28[21], tmp28[20], tmp28[19], tmp28[18], tmp28[17], tmp28[16], tmp28[15], tmp28[14], tmp28[13], tmp28[12], tmp28[11], tmp28[10], tmp28[9], tmp28[8], tmp28[7], tmp28[6], tmp28[5], tmp28[4], tmp28[3], tmp28[2], tmp28[1]};
    assign tmp2885 = {tmp2884[254]};
    assign tmp2886 = {tmp2885};
    assign tmp2887 = {tmp2886, tmp2884};
    assign tmp2888 = ~tmp35;
    assign tmp2889 = ~tmp36;
    assign tmp2890 = tmp2888 & tmp2889;
    assign tmp2891 = ~tmp57;
    assign tmp2892 = tmp2890 & tmp2891;
    assign tmp2893 = ~tmp1034;
    assign tmp2894 = tmp2892 & tmp2893;
    assign tmp2895 = tmp2894 & tmp2071;
    assign tmp2896 = ~tmp2583;
    assign tmp2897 = tmp2895 & tmp2896;
    assign tmp2898 = tmp2897 & tmp23;
    assign tmp2899 = ~tmp2627;
    assign tmp2900 = tmp2898 & tmp2899;
    assign tmp2901 = tmp2900 & tmp2798;
    assign tmp2902 = tmp2901 & tmp24;
    assign tmp2903 = ~tmp35;
    assign tmp2904 = ~tmp36;
    assign tmp2905 = tmp2903 & tmp2904;
    assign tmp2906 = ~tmp57;
    assign tmp2907 = tmp2905 & tmp2906;
    assign tmp2908 = ~tmp1034;
    assign tmp2909 = tmp2907 & tmp2908;
    assign tmp2910 = tmp2909 & tmp2071;
    assign tmp2911 = ~tmp2583;
    assign tmp2912 = tmp2910 & tmp2911;
    assign tmp2913 = tmp2912 & tmp23;
    assign tmp2914 = ~tmp2627;
    assign tmp2915 = tmp2913 & tmp2914;
    assign tmp2916 = tmp2915 & tmp2798;
    assign tmp2917 = tmp2916 & tmp24;
    assign tmp2918 = ~tmp35;
    assign tmp2919 = ~tmp36;
    assign tmp2920 = tmp2918 & tmp2919;
    assign tmp2921 = ~tmp57;
    assign tmp2922 = tmp2920 & tmp2921;
    assign tmp2923 = ~tmp1034;
    assign tmp2924 = tmp2922 & tmp2923;
    assign tmp2925 = tmp2924 & tmp2071;
    assign tmp2926 = ~tmp2583;
    assign tmp2927 = tmp2925 & tmp2926;
    assign tmp2928 = tmp2927 & tmp23;
    assign tmp2929 = ~tmp2627;
    assign tmp2930 = tmp2928 & tmp2929;
    assign tmp2931 = tmp2930 & tmp2798;
    assign tmp2932 = tmp2931 & tmp24;
    assign tmp2933 = ~tmp35;
    assign tmp2934 = ~tmp36;
    assign tmp2935 = tmp2933 & tmp2934;
    assign tmp2936 = ~tmp57;
    assign tmp2937 = tmp2935 & tmp2936;
    assign tmp2938 = ~tmp1034;
    assign tmp2939 = tmp2937 & tmp2938;
    assign tmp2940 = tmp2939 & tmp2071;
    assign tmp2941 = ~tmp2583;
    assign tmp2942 = tmp2940 & tmp2941;
    assign tmp2943 = tmp2942 & tmp23;
    assign tmp2944 = ~tmp2627;
    assign tmp2945 = tmp2943 & tmp2944;
    assign tmp2946 = tmp2945 & tmp2798;
    assign tmp2947 = tmp2946 & tmp24;
    assign tmp2948 = ~tmp35;
    assign tmp2949 = ~tmp36;
    assign tmp2950 = tmp2948 & tmp2949;
    assign tmp2951 = ~tmp57;
    assign tmp2952 = tmp2950 & tmp2951;
    assign tmp2953 = ~tmp1034;
    assign tmp2954 = tmp2952 & tmp2953;
    assign tmp2955 = tmp2954 & tmp2071;
    assign tmp2956 = ~tmp2583;
    assign tmp2957 = tmp2955 & tmp2956;
    assign tmp2958 = tmp2957 & tmp23;
    assign tmp2959 = ~tmp2627;
    assign tmp2960 = tmp2958 & tmp2959;
    assign tmp2961 = tmp2960 & tmp2798;
    assign tmp2962 = tmp2961 & tmp24;
    assign tmp2963 = ~tmp35;
    assign tmp2964 = ~tmp36;
    assign tmp2965 = tmp2963 & tmp2964;
    assign tmp2966 = ~tmp57;
    assign tmp2967 = tmp2965 & tmp2966;
    assign tmp2968 = ~tmp1034;
    assign tmp2969 = tmp2967 & tmp2968;
    assign tmp2970 = tmp2969 & tmp2071;
    assign tmp2971 = ~tmp2583;
    assign tmp2972 = tmp2970 & tmp2971;
    assign tmp2973 = tmp2972 & tmp23;
    assign tmp2974 = ~tmp2627;
    assign tmp2975 = tmp2973 & tmp2974;
    assign tmp2976 = tmp2975 & tmp2798;
    assign tmp2977 = ~tmp24;
    assign tmp2978 = tmp2976 & tmp2977;
    assign tmp2979 = ~tmp35;
    assign tmp2980 = ~tmp36;
    assign tmp2981 = tmp2979 & tmp2980;
    assign tmp2982 = ~tmp57;
    assign tmp2983 = tmp2981 & tmp2982;
    assign tmp2984 = ~tmp1034;
    assign tmp2985 = tmp2983 & tmp2984;
    assign tmp2986 = tmp2985 & tmp2071;
    assign tmp2987 = ~tmp2583;
    assign tmp2988 = tmp2986 & tmp2987;
    assign tmp2989 = tmp2988 & tmp23;
    assign tmp2990 = ~tmp2627;
    assign tmp2991 = tmp2989 & tmp2990;
    assign tmp2992 = tmp2991 & tmp2798;
    assign tmp2993 = ~tmp24;
    assign tmp2994 = tmp2992 & tmp2993;
    assign tmp2995 = ~tmp35;
    assign tmp2996 = ~tmp36;
    assign tmp2997 = tmp2995 & tmp2996;
    assign tmp2998 = ~tmp57;
    assign tmp2999 = tmp2997 & tmp2998;
    assign tmp3000 = ~tmp1034;
    assign tmp3001 = tmp2999 & tmp3000;
    assign tmp3002 = tmp3001 & tmp2071;
    assign tmp3003 = ~tmp2583;
    assign tmp3004 = tmp3002 & tmp3003;
    assign tmp3005 = tmp3004 & tmp23;
    assign tmp3006 = ~tmp2627;
    assign tmp3007 = tmp3005 & tmp3006;
    assign tmp3008 = tmp3007 & tmp2798;
    assign tmp3009 = ~tmp24;
    assign tmp3010 = tmp3008 & tmp3009;
    assign tmp3011 = ~tmp35;
    assign tmp3012 = ~tmp36;
    assign tmp3013 = tmp3011 & tmp3012;
    assign tmp3014 = ~tmp57;
    assign tmp3015 = tmp3013 & tmp3014;
    assign tmp3016 = ~tmp1034;
    assign tmp3017 = tmp3015 & tmp3016;
    assign tmp3018 = tmp3017 & tmp2071;
    assign tmp3019 = ~tmp2583;
    assign tmp3020 = tmp3018 & tmp3019;
    assign tmp3021 = tmp3020 & tmp23;
    assign tmp3022 = ~tmp2627;
    assign tmp3023 = tmp3021 & tmp3022;
    assign tmp3024 = tmp3023 & tmp2798;
    assign tmp3025 = ~tmp24;
    assign tmp3026 = tmp3024 & tmp3025;
    assign tmp3027 = {tmp29[254], tmp29[253], tmp29[252], tmp29[251], tmp29[250], tmp29[249], tmp29[248], tmp29[247], tmp29[246], tmp29[245], tmp29[244], tmp29[243], tmp29[242], tmp29[241], tmp29[240], tmp29[239], tmp29[238], tmp29[237], tmp29[236], tmp29[235], tmp29[234], tmp29[233], tmp29[232], tmp29[231], tmp29[230], tmp29[229], tmp29[228], tmp29[227], tmp29[226], tmp29[225], tmp29[224], tmp29[223], tmp29[222], tmp29[221], tmp29[220], tmp29[219], tmp29[218], tmp29[217], tmp29[216], tmp29[215], tmp29[214], tmp29[213], tmp29[212], tmp29[211], tmp29[210], tmp29[209], tmp29[208], tmp29[207], tmp29[206], tmp29[205], tmp29[204], tmp29[203], tmp29[202], tmp29[201], tmp29[200], tmp29[199], tmp29[198], tmp29[197], tmp29[196], tmp29[195], tmp29[194], tmp29[193], tmp29[192], tmp29[191], tmp29[190], tmp29[189], tmp29[188], tmp29[187], tmp29[186], tmp29[185], tmp29[184], tmp29[183], tmp29[182], tmp29[181], tmp29[180], tmp29[179], tmp29[178], tmp29[177], tmp29[176], tmp29[175], tmp29[174], tmp29[173], tmp29[172], tmp29[171], tmp29[170], tmp29[169], tmp29[168], tmp29[167], tmp29[166], tmp29[165], tmp29[164], tmp29[163], tmp29[162], tmp29[161], tmp29[160], tmp29[159], tmp29[158], tmp29[157], tmp29[156], tmp29[155], tmp29[154], tmp29[153], tmp29[152], tmp29[151], tmp29[150], tmp29[149], tmp29[148], tmp29[147], tmp29[146], tmp29[145], tmp29[144], tmp29[143], tmp29[142], tmp29[141], tmp29[140], tmp29[139], tmp29[138], tmp29[137], tmp29[136], tmp29[135], tmp29[134], tmp29[133], tmp29[132], tmp29[131], tmp29[130], tmp29[129], tmp29[128], tmp29[127], tmp29[126], tmp29[125], tmp29[124], tmp29[123], tmp29[122], tmp29[121], tmp29[120], tmp29[119], tmp29[118], tmp29[117], tmp29[116], tmp29[115], tmp29[114], tmp29[113], tmp29[112], tmp29[111], tmp29[110], tmp29[109], tmp29[108], tmp29[107], tmp29[106], tmp29[105], tmp29[104], tmp29[103], tmp29[102], tmp29[101], tmp29[100], tmp29[99], tmp29[98], tmp29[97], tmp29[96], tmp29[95], tmp29[94], tmp29[93], tmp29[92], tmp29[91], tmp29[90], tmp29[89], tmp29[88], tmp29[87], tmp29[86], tmp29[85], tmp29[84], tmp29[83], tmp29[82], tmp29[81], tmp29[80], tmp29[79], tmp29[78], tmp29[77], tmp29[76], tmp29[75], tmp29[74], tmp29[73], tmp29[72], tmp29[71], tmp29[70], tmp29[69], tmp29[68], tmp29[67], tmp29[66], tmp29[65], tmp29[64], tmp29[63], tmp29[62], tmp29[61], tmp29[60], tmp29[59], tmp29[58], tmp29[57], tmp29[56], tmp29[55], tmp29[54], tmp29[53], tmp29[52], tmp29[51], tmp29[50], tmp29[49], tmp29[48], tmp29[47], tmp29[46], tmp29[45], tmp29[44], tmp29[43], tmp29[42], tmp29[41], tmp29[40], tmp29[39], tmp29[38], tmp29[37], tmp29[36], tmp29[35], tmp29[34], tmp29[33], tmp29[32], tmp29[31], tmp29[30], tmp29[29], tmp29[28], tmp29[27], tmp29[26], tmp29[25], tmp29[24], tmp29[23], tmp29[22], tmp29[21], tmp29[20], tmp29[19], tmp29[18], tmp29[17], tmp29[16], tmp29[15], tmp29[14], tmp29[13], tmp29[12], tmp29[11], tmp29[10], tmp29[9], tmp29[8], tmp29[7], tmp29[6], tmp29[5], tmp29[4], tmp29[3], tmp29[2], tmp29[1], tmp29[0]};
    assign tmp3028 = {tmp3027, const_319_0};
    assign tmp3029 = {const_320_0};
    assign tmp3030 = {tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029, tmp3029};
    assign tmp3031 = {tmp3030, const_320_0};
    assign tmp3032 = {tmp29[255]};
    assign tmp3033 = tmp3031 - tmp29;
    assign tmp3034 = {tmp3033[256]};
    assign tmp3035 = {tmp3031[255]};
    assign tmp3036 = ~tmp3035;
    assign tmp3037 = tmp3034 ^ tmp3036;
    assign tmp3038 = {tmp29[255]};
    assign tmp3039 = ~tmp3038;
    assign tmp3040 = tmp3037 ^ tmp3039;
    assign tmp3041 = {tmp3028[255]};
    assign tmp3042 = {const_321_0};
    assign tmp3043 = {tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042, tmp3042};
    assign tmp3044 = {tmp3043, const_321_0};
    assign tmp3045 = tmp3028 - tmp3044;
    assign tmp3046 = {tmp3045[256]};
    assign tmp3047 = {tmp3028[255]};
    assign tmp3048 = ~tmp3047;
    assign tmp3049 = tmp3046 ^ tmp3048;
    assign tmp3050 = {tmp3044[255]};
    assign tmp3051 = ~tmp3050;
    assign tmp3052 = tmp3049 ^ tmp3051;
    assign tmp3053 = tmp3040 & tmp3052;
    assign tmp3054 = {tmp29[255]};
    assign tmp3055 = {const_322_0};
    assign tmp3056 = {tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055, tmp3055};
    assign tmp3057 = {tmp3056, const_322_0};
    assign tmp3058 = tmp29 - tmp3057;
    assign tmp3059 = {tmp3058[256]};
    assign tmp3060 = {tmp29[255]};
    assign tmp3061 = ~tmp3060;
    assign tmp3062 = tmp3059 ^ tmp3061;
    assign tmp3063 = {tmp3057[255]};
    assign tmp3064 = ~tmp3063;
    assign tmp3065 = tmp3062 ^ tmp3064;
    assign tmp3066 = {const_323_0};
    assign tmp3067 = {tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066, tmp3066};
    assign tmp3068 = {tmp3067, const_323_0};
    assign tmp3069 = {tmp3028[255]};
    assign tmp3070 = tmp3068 - tmp3028;
    assign tmp3071 = {tmp3070[256]};
    assign tmp3072 = {tmp3068[255]};
    assign tmp3073 = ~tmp3072;
    assign tmp3074 = tmp3071 ^ tmp3073;
    assign tmp3075 = {tmp3028[255]};
    assign tmp3076 = ~tmp3075;
    assign tmp3077 = tmp3074 ^ tmp3076;
    assign tmp3078 = tmp3068 == tmp3028;
    assign tmp3079 = tmp3077 | tmp3078;
    assign tmp3080 = tmp3065 & tmp3079;
    assign tmp3081 = tmp3053 ? const_324_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp3028;
    assign tmp3082 = tmp3080 ? _ver_out_tmp_23 : tmp3081;
    assign tmp3083 = ~tmp35;
    assign tmp3084 = ~tmp36;
    assign tmp3085 = tmp3083 & tmp3084;
    assign tmp3086 = ~tmp57;
    assign tmp3087 = tmp3085 & tmp3086;
    assign tmp3088 = ~tmp1034;
    assign tmp3089 = tmp3087 & tmp3088;
    assign tmp3090 = tmp3089 & tmp2071;
    assign tmp3091 = ~tmp2583;
    assign tmp3092 = tmp3090 & tmp3091;
    assign tmp3093 = tmp3092 & tmp23;
    assign tmp3094 = ~tmp2627;
    assign tmp3095 = tmp3093 & tmp3094;
    assign tmp3096 = tmp3095 & tmp2798;
    assign tmp3097 = ~tmp24;
    assign tmp3098 = tmp3096 & tmp3097;
    assign tmp3099 = {tmp30[254], tmp30[253], tmp30[252], tmp30[251], tmp30[250], tmp30[249], tmp30[248], tmp30[247], tmp30[246], tmp30[245], tmp30[244], tmp30[243], tmp30[242], tmp30[241], tmp30[240], tmp30[239], tmp30[238], tmp30[237], tmp30[236], tmp30[235], tmp30[234], tmp30[233], tmp30[232], tmp30[231], tmp30[230], tmp30[229], tmp30[228], tmp30[227], tmp30[226], tmp30[225], tmp30[224], tmp30[223], tmp30[222], tmp30[221], tmp30[220], tmp30[219], tmp30[218], tmp30[217], tmp30[216], tmp30[215], tmp30[214], tmp30[213], tmp30[212], tmp30[211], tmp30[210], tmp30[209], tmp30[208], tmp30[207], tmp30[206], tmp30[205], tmp30[204], tmp30[203], tmp30[202], tmp30[201], tmp30[200], tmp30[199], tmp30[198], tmp30[197], tmp30[196], tmp30[195], tmp30[194], tmp30[193], tmp30[192], tmp30[191], tmp30[190], tmp30[189], tmp30[188], tmp30[187], tmp30[186], tmp30[185], tmp30[184], tmp30[183], tmp30[182], tmp30[181], tmp30[180], tmp30[179], tmp30[178], tmp30[177], tmp30[176], tmp30[175], tmp30[174], tmp30[173], tmp30[172], tmp30[171], tmp30[170], tmp30[169], tmp30[168], tmp30[167], tmp30[166], tmp30[165], tmp30[164], tmp30[163], tmp30[162], tmp30[161], tmp30[160], tmp30[159], tmp30[158], tmp30[157], tmp30[156], tmp30[155], tmp30[154], tmp30[153], tmp30[152], tmp30[151], tmp30[150], tmp30[149], tmp30[148], tmp30[147], tmp30[146], tmp30[145], tmp30[144], tmp30[143], tmp30[142], tmp30[141], tmp30[140], tmp30[139], tmp30[138], tmp30[137], tmp30[136], tmp30[135], tmp30[134], tmp30[133], tmp30[132], tmp30[131], tmp30[130], tmp30[129], tmp30[128], tmp30[127], tmp30[126], tmp30[125], tmp30[124], tmp30[123], tmp30[122], tmp30[121], tmp30[120], tmp30[119], tmp30[118], tmp30[117], tmp30[116], tmp30[115], tmp30[114], tmp30[113], tmp30[112], tmp30[111], tmp30[110], tmp30[109], tmp30[108], tmp30[107], tmp30[106], tmp30[105], tmp30[104], tmp30[103], tmp30[102], tmp30[101], tmp30[100], tmp30[99], tmp30[98], tmp30[97], tmp30[96], tmp30[95], tmp30[94], tmp30[93], tmp30[92], tmp30[91], tmp30[90], tmp30[89], tmp30[88], tmp30[87], tmp30[86], tmp30[85], tmp30[84], tmp30[83], tmp30[82], tmp30[81], tmp30[80], tmp30[79], tmp30[78], tmp30[77], tmp30[76], tmp30[75], tmp30[74], tmp30[73], tmp30[72], tmp30[71], tmp30[70], tmp30[69], tmp30[68], tmp30[67], tmp30[66], tmp30[65], tmp30[64], tmp30[63], tmp30[62], tmp30[61], tmp30[60], tmp30[59], tmp30[58], tmp30[57], tmp30[56], tmp30[55], tmp30[54], tmp30[53], tmp30[52], tmp30[51], tmp30[50], tmp30[49], tmp30[48], tmp30[47], tmp30[46], tmp30[45], tmp30[44], tmp30[43], tmp30[42], tmp30[41], tmp30[40], tmp30[39], tmp30[38], tmp30[37], tmp30[36], tmp30[35], tmp30[34], tmp30[33], tmp30[32], tmp30[31], tmp30[30], tmp30[29], tmp30[28], tmp30[27], tmp30[26], tmp30[25], tmp30[24], tmp30[23], tmp30[22], tmp30[21], tmp30[20], tmp30[19], tmp30[18], tmp30[17], tmp30[16], tmp30[15], tmp30[14], tmp30[13], tmp30[12], tmp30[11], tmp30[10], tmp30[9], tmp30[8], tmp30[7], tmp30[6], tmp30[5], tmp30[4], tmp30[3], tmp30[2], tmp30[1], tmp30[0]};
    assign tmp3100 = {tmp3099, const_326_0};
    assign tmp3101 = {const_327_0};
    assign tmp3102 = {tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101, tmp3101};
    assign tmp3103 = {tmp3102, const_327_0};
    assign tmp3104 = {tmp30[255]};
    assign tmp3105 = tmp3103 - tmp30;
    assign tmp3106 = {tmp3105[256]};
    assign tmp3107 = {tmp3103[255]};
    assign tmp3108 = ~tmp3107;
    assign tmp3109 = tmp3106 ^ tmp3108;
    assign tmp3110 = {tmp30[255]};
    assign tmp3111 = ~tmp3110;
    assign tmp3112 = tmp3109 ^ tmp3111;
    assign tmp3113 = {tmp3100[255]};
    assign tmp3114 = {const_328_0};
    assign tmp3115 = {tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114, tmp3114};
    assign tmp3116 = {tmp3115, const_328_0};
    assign tmp3117 = tmp3100 - tmp3116;
    assign tmp3118 = {tmp3117[256]};
    assign tmp3119 = {tmp3100[255]};
    assign tmp3120 = ~tmp3119;
    assign tmp3121 = tmp3118 ^ tmp3120;
    assign tmp3122 = {tmp3116[255]};
    assign tmp3123 = ~tmp3122;
    assign tmp3124 = tmp3121 ^ tmp3123;
    assign tmp3125 = tmp3112 & tmp3124;
    assign tmp3126 = {tmp30[255]};
    assign tmp3127 = {const_329_0};
    assign tmp3128 = {tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127, tmp3127};
    assign tmp3129 = {tmp3128, const_329_0};
    assign tmp3130 = tmp30 - tmp3129;
    assign tmp3131 = {tmp3130[256]};
    assign tmp3132 = {tmp30[255]};
    assign tmp3133 = ~tmp3132;
    assign tmp3134 = tmp3131 ^ tmp3133;
    assign tmp3135 = {tmp3129[255]};
    assign tmp3136 = ~tmp3135;
    assign tmp3137 = tmp3134 ^ tmp3136;
    assign tmp3138 = {const_330_0};
    assign tmp3139 = {tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138, tmp3138};
    assign tmp3140 = {tmp3139, const_330_0};
    assign tmp3141 = {tmp3100[255]};
    assign tmp3142 = tmp3140 - tmp3100;
    assign tmp3143 = {tmp3142[256]};
    assign tmp3144 = {tmp3140[255]};
    assign tmp3145 = ~tmp3144;
    assign tmp3146 = tmp3143 ^ tmp3145;
    assign tmp3147 = {tmp3100[255]};
    assign tmp3148 = ~tmp3147;
    assign tmp3149 = tmp3146 ^ tmp3148;
    assign tmp3150 = tmp3140 == tmp3100;
    assign tmp3151 = tmp3149 | tmp3150;
    assign tmp3152 = tmp3137 & tmp3151;
    assign tmp3153 = tmp3125 ? const_331_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp3100;
    assign tmp3154 = tmp3152 ? _ver_out_tmp_71 : tmp3153;
    assign tmp3155 = ~tmp35;
    assign tmp3156 = ~tmp36;
    assign tmp3157 = tmp3155 & tmp3156;
    assign tmp3158 = ~tmp57;
    assign tmp3159 = tmp3157 & tmp3158;
    assign tmp3160 = ~tmp1034;
    assign tmp3161 = tmp3159 & tmp3160;
    assign tmp3162 = tmp3161 & tmp2071;
    assign tmp3163 = ~tmp2583;
    assign tmp3164 = tmp3162 & tmp3163;
    assign tmp3165 = tmp3164 & tmp23;
    assign tmp3166 = ~tmp2627;
    assign tmp3167 = tmp3165 & tmp3166;
    assign tmp3168 = tmp3167 & tmp2798;
    assign tmp3169 = ~tmp24;
    assign tmp3170 = tmp3168 & tmp3169;
    assign tmp3171 = {tmp31[254], tmp31[253], tmp31[252], tmp31[251], tmp31[250], tmp31[249], tmp31[248], tmp31[247], tmp31[246], tmp31[245], tmp31[244], tmp31[243], tmp31[242], tmp31[241], tmp31[240], tmp31[239], tmp31[238], tmp31[237], tmp31[236], tmp31[235], tmp31[234], tmp31[233], tmp31[232], tmp31[231], tmp31[230], tmp31[229], tmp31[228], tmp31[227], tmp31[226], tmp31[225], tmp31[224], tmp31[223], tmp31[222], tmp31[221], tmp31[220], tmp31[219], tmp31[218], tmp31[217], tmp31[216], tmp31[215], tmp31[214], tmp31[213], tmp31[212], tmp31[211], tmp31[210], tmp31[209], tmp31[208], tmp31[207], tmp31[206], tmp31[205], tmp31[204], tmp31[203], tmp31[202], tmp31[201], tmp31[200], tmp31[199], tmp31[198], tmp31[197], tmp31[196], tmp31[195], tmp31[194], tmp31[193], tmp31[192], tmp31[191], tmp31[190], tmp31[189], tmp31[188], tmp31[187], tmp31[186], tmp31[185], tmp31[184], tmp31[183], tmp31[182], tmp31[181], tmp31[180], tmp31[179], tmp31[178], tmp31[177], tmp31[176], tmp31[175], tmp31[174], tmp31[173], tmp31[172], tmp31[171], tmp31[170], tmp31[169], tmp31[168], tmp31[167], tmp31[166], tmp31[165], tmp31[164], tmp31[163], tmp31[162], tmp31[161], tmp31[160], tmp31[159], tmp31[158], tmp31[157], tmp31[156], tmp31[155], tmp31[154], tmp31[153], tmp31[152], tmp31[151], tmp31[150], tmp31[149], tmp31[148], tmp31[147], tmp31[146], tmp31[145], tmp31[144], tmp31[143], tmp31[142], tmp31[141], tmp31[140], tmp31[139], tmp31[138], tmp31[137], tmp31[136], tmp31[135], tmp31[134], tmp31[133], tmp31[132], tmp31[131], tmp31[130], tmp31[129], tmp31[128], tmp31[127], tmp31[126], tmp31[125], tmp31[124], tmp31[123], tmp31[122], tmp31[121], tmp31[120], tmp31[119], tmp31[118], tmp31[117], tmp31[116], tmp31[115], tmp31[114], tmp31[113], tmp31[112], tmp31[111], tmp31[110], tmp31[109], tmp31[108], tmp31[107], tmp31[106], tmp31[105], tmp31[104], tmp31[103], tmp31[102], tmp31[101], tmp31[100], tmp31[99], tmp31[98], tmp31[97], tmp31[96], tmp31[95], tmp31[94], tmp31[93], tmp31[92], tmp31[91], tmp31[90], tmp31[89], tmp31[88], tmp31[87], tmp31[86], tmp31[85], tmp31[84], tmp31[83], tmp31[82], tmp31[81], tmp31[80], tmp31[79], tmp31[78], tmp31[77], tmp31[76], tmp31[75], tmp31[74], tmp31[73], tmp31[72], tmp31[71], tmp31[70], tmp31[69], tmp31[68], tmp31[67], tmp31[66], tmp31[65], tmp31[64], tmp31[63], tmp31[62], tmp31[61], tmp31[60], tmp31[59], tmp31[58], tmp31[57], tmp31[56], tmp31[55], tmp31[54], tmp31[53], tmp31[52], tmp31[51], tmp31[50], tmp31[49], tmp31[48], tmp31[47], tmp31[46], tmp31[45], tmp31[44], tmp31[43], tmp31[42], tmp31[41], tmp31[40], tmp31[39], tmp31[38], tmp31[37], tmp31[36], tmp31[35], tmp31[34], tmp31[33], tmp31[32], tmp31[31], tmp31[30], tmp31[29], tmp31[28], tmp31[27], tmp31[26], tmp31[25], tmp31[24], tmp31[23], tmp31[22], tmp31[21], tmp31[20], tmp31[19], tmp31[18], tmp31[17], tmp31[16], tmp31[15], tmp31[14], tmp31[13], tmp31[12], tmp31[11], tmp31[10], tmp31[9], tmp31[8], tmp31[7], tmp31[6], tmp31[5], tmp31[4], tmp31[3], tmp31[2], tmp31[1], tmp31[0]};
    assign tmp3172 = {tmp3171, const_333_0};
    assign tmp3173 = {const_334_0};
    assign tmp3174 = {tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173, tmp3173};
    assign tmp3175 = {tmp3174, const_334_0};
    assign tmp3176 = {tmp31[255]};
    assign tmp3177 = tmp3175 - tmp31;
    assign tmp3178 = {tmp3177[256]};
    assign tmp3179 = {tmp3175[255]};
    assign tmp3180 = ~tmp3179;
    assign tmp3181 = tmp3178 ^ tmp3180;
    assign tmp3182 = {tmp31[255]};
    assign tmp3183 = ~tmp3182;
    assign tmp3184 = tmp3181 ^ tmp3183;
    assign tmp3185 = {tmp3172[255]};
    assign tmp3186 = {const_335_0};
    assign tmp3187 = {tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186, tmp3186};
    assign tmp3188 = {tmp3187, const_335_0};
    assign tmp3189 = tmp3172 - tmp3188;
    assign tmp3190 = {tmp3189[256]};
    assign tmp3191 = {tmp3172[255]};
    assign tmp3192 = ~tmp3191;
    assign tmp3193 = tmp3190 ^ tmp3192;
    assign tmp3194 = {tmp3188[255]};
    assign tmp3195 = ~tmp3194;
    assign tmp3196 = tmp3193 ^ tmp3195;
    assign tmp3197 = tmp3184 & tmp3196;
    assign tmp3198 = {tmp31[255]};
    assign tmp3199 = {const_336_0};
    assign tmp3200 = {tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199, tmp3199};
    assign tmp3201 = {tmp3200, const_336_0};
    assign tmp3202 = tmp31 - tmp3201;
    assign tmp3203 = {tmp3202[256]};
    assign tmp3204 = {tmp31[255]};
    assign tmp3205 = ~tmp3204;
    assign tmp3206 = tmp3203 ^ tmp3205;
    assign tmp3207 = {tmp3201[255]};
    assign tmp3208 = ~tmp3207;
    assign tmp3209 = tmp3206 ^ tmp3208;
    assign tmp3210 = {const_337_0};
    assign tmp3211 = {tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210, tmp3210};
    assign tmp3212 = {tmp3211, const_337_0};
    assign tmp3213 = {tmp3172[255]};
    assign tmp3214 = tmp3212 - tmp3172;
    assign tmp3215 = {tmp3214[256]};
    assign tmp3216 = {tmp3212[255]};
    assign tmp3217 = ~tmp3216;
    assign tmp3218 = tmp3215 ^ tmp3217;
    assign tmp3219 = {tmp3172[255]};
    assign tmp3220 = ~tmp3219;
    assign tmp3221 = tmp3218 ^ tmp3220;
    assign tmp3222 = tmp3212 == tmp3172;
    assign tmp3223 = tmp3221 | tmp3222;
    assign tmp3224 = tmp3209 & tmp3223;
    assign tmp3225 = tmp3197 ? const_338_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp3172;
    assign tmp3226 = tmp3224 ? _ver_out_tmp_72 : tmp3225;
    assign tmp3227 = ~tmp35;
    assign tmp3228 = ~tmp36;
    assign tmp3229 = tmp3227 & tmp3228;
    assign tmp3230 = ~tmp57;
    assign tmp3231 = tmp3229 & tmp3230;
    assign tmp3232 = ~tmp1034;
    assign tmp3233 = tmp3231 & tmp3232;
    assign tmp3234 = tmp3233 & tmp2071;
    assign tmp3235 = ~tmp2583;
    assign tmp3236 = tmp3234 & tmp3235;
    assign tmp3237 = tmp3236 & tmp23;
    assign tmp3238 = ~tmp2627;
    assign tmp3239 = tmp3237 & tmp3238;
    assign tmp3240 = tmp3239 & tmp2798;
    assign tmp3241 = ~tmp24;
    assign tmp3242 = tmp3240 & tmp3241;
    assign tmp3243 = {tmp32[254], tmp32[253], tmp32[252], tmp32[251], tmp32[250], tmp32[249], tmp32[248], tmp32[247], tmp32[246], tmp32[245], tmp32[244], tmp32[243], tmp32[242], tmp32[241], tmp32[240], tmp32[239], tmp32[238], tmp32[237], tmp32[236], tmp32[235], tmp32[234], tmp32[233], tmp32[232], tmp32[231], tmp32[230], tmp32[229], tmp32[228], tmp32[227], tmp32[226], tmp32[225], tmp32[224], tmp32[223], tmp32[222], tmp32[221], tmp32[220], tmp32[219], tmp32[218], tmp32[217], tmp32[216], tmp32[215], tmp32[214], tmp32[213], tmp32[212], tmp32[211], tmp32[210], tmp32[209], tmp32[208], tmp32[207], tmp32[206], tmp32[205], tmp32[204], tmp32[203], tmp32[202], tmp32[201], tmp32[200], tmp32[199], tmp32[198], tmp32[197], tmp32[196], tmp32[195], tmp32[194], tmp32[193], tmp32[192], tmp32[191], tmp32[190], tmp32[189], tmp32[188], tmp32[187], tmp32[186], tmp32[185], tmp32[184], tmp32[183], tmp32[182], tmp32[181], tmp32[180], tmp32[179], tmp32[178], tmp32[177], tmp32[176], tmp32[175], tmp32[174], tmp32[173], tmp32[172], tmp32[171], tmp32[170], tmp32[169], tmp32[168], tmp32[167], tmp32[166], tmp32[165], tmp32[164], tmp32[163], tmp32[162], tmp32[161], tmp32[160], tmp32[159], tmp32[158], tmp32[157], tmp32[156], tmp32[155], tmp32[154], tmp32[153], tmp32[152], tmp32[151], tmp32[150], tmp32[149], tmp32[148], tmp32[147], tmp32[146], tmp32[145], tmp32[144], tmp32[143], tmp32[142], tmp32[141], tmp32[140], tmp32[139], tmp32[138], tmp32[137], tmp32[136], tmp32[135], tmp32[134], tmp32[133], tmp32[132], tmp32[131], tmp32[130], tmp32[129], tmp32[128], tmp32[127], tmp32[126], tmp32[125], tmp32[124], tmp32[123], tmp32[122], tmp32[121], tmp32[120], tmp32[119], tmp32[118], tmp32[117], tmp32[116], tmp32[115], tmp32[114], tmp32[113], tmp32[112], tmp32[111], tmp32[110], tmp32[109], tmp32[108], tmp32[107], tmp32[106], tmp32[105], tmp32[104], tmp32[103], tmp32[102], tmp32[101], tmp32[100], tmp32[99], tmp32[98], tmp32[97], tmp32[96], tmp32[95], tmp32[94], tmp32[93], tmp32[92], tmp32[91], tmp32[90], tmp32[89], tmp32[88], tmp32[87], tmp32[86], tmp32[85], tmp32[84], tmp32[83], tmp32[82], tmp32[81], tmp32[80], tmp32[79], tmp32[78], tmp32[77], tmp32[76], tmp32[75], tmp32[74], tmp32[73], tmp32[72], tmp32[71], tmp32[70], tmp32[69], tmp32[68], tmp32[67], tmp32[66], tmp32[65], tmp32[64], tmp32[63], tmp32[62], tmp32[61], tmp32[60], tmp32[59], tmp32[58], tmp32[57], tmp32[56], tmp32[55], tmp32[54], tmp32[53], tmp32[52], tmp32[51], tmp32[50], tmp32[49], tmp32[48], tmp32[47], tmp32[46], tmp32[45], tmp32[44], tmp32[43], tmp32[42], tmp32[41], tmp32[40], tmp32[39], tmp32[38], tmp32[37], tmp32[36], tmp32[35], tmp32[34], tmp32[33], tmp32[32], tmp32[31], tmp32[30], tmp32[29], tmp32[28], tmp32[27], tmp32[26], tmp32[25], tmp32[24], tmp32[23], tmp32[22], tmp32[21], tmp32[20], tmp32[19], tmp32[18], tmp32[17], tmp32[16], tmp32[15], tmp32[14], tmp32[13], tmp32[12], tmp32[11], tmp32[10], tmp32[9], tmp32[8], tmp32[7], tmp32[6], tmp32[5], tmp32[4], tmp32[3], tmp32[2], tmp32[1], tmp32[0]};
    assign tmp3244 = {tmp3243, const_340_0};
    assign tmp3245 = {const_341_0};
    assign tmp3246 = {tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245, tmp3245};
    assign tmp3247 = {tmp3246, const_341_0};
    assign tmp3248 = {tmp32[255]};
    assign tmp3249 = tmp3247 - tmp32;
    assign tmp3250 = {tmp3249[256]};
    assign tmp3251 = {tmp3247[255]};
    assign tmp3252 = ~tmp3251;
    assign tmp3253 = tmp3250 ^ tmp3252;
    assign tmp3254 = {tmp32[255]};
    assign tmp3255 = ~tmp3254;
    assign tmp3256 = tmp3253 ^ tmp3255;
    assign tmp3257 = {tmp3244[255]};
    assign tmp3258 = {const_342_0};
    assign tmp3259 = {tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258, tmp3258};
    assign tmp3260 = {tmp3259, const_342_0};
    assign tmp3261 = tmp3244 - tmp3260;
    assign tmp3262 = {tmp3261[256]};
    assign tmp3263 = {tmp3244[255]};
    assign tmp3264 = ~tmp3263;
    assign tmp3265 = tmp3262 ^ tmp3264;
    assign tmp3266 = {tmp3260[255]};
    assign tmp3267 = ~tmp3266;
    assign tmp3268 = tmp3265 ^ tmp3267;
    assign tmp3269 = tmp3256 & tmp3268;
    assign tmp3270 = {tmp32[255]};
    assign tmp3271 = {const_343_0};
    assign tmp3272 = {tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271, tmp3271};
    assign tmp3273 = {tmp3272, const_343_0};
    assign tmp3274 = tmp32 - tmp3273;
    assign tmp3275 = {tmp3274[256]};
    assign tmp3276 = {tmp32[255]};
    assign tmp3277 = ~tmp3276;
    assign tmp3278 = tmp3275 ^ tmp3277;
    assign tmp3279 = {tmp3273[255]};
    assign tmp3280 = ~tmp3279;
    assign tmp3281 = tmp3278 ^ tmp3280;
    assign tmp3282 = {const_344_0};
    assign tmp3283 = {tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282, tmp3282};
    assign tmp3284 = {tmp3283, const_344_0};
    assign tmp3285 = {tmp3244[255]};
    assign tmp3286 = tmp3284 - tmp3244;
    assign tmp3287 = {tmp3286[256]};
    assign tmp3288 = {tmp3284[255]};
    assign tmp3289 = ~tmp3288;
    assign tmp3290 = tmp3287 ^ tmp3289;
    assign tmp3291 = {tmp3244[255]};
    assign tmp3292 = ~tmp3291;
    assign tmp3293 = tmp3290 ^ tmp3292;
    assign tmp3294 = tmp3284 == tmp3244;
    assign tmp3295 = tmp3293 | tmp3294;
    assign tmp3296 = tmp3281 & tmp3295;
    assign tmp3297 = tmp3269 ? const_345_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp3244;
    assign tmp3298 = tmp3296 ? _ver_out_tmp_75 : tmp3297;
    assign tmp3299 = ~tmp35;
    assign tmp3300 = ~tmp36;
    assign tmp3301 = tmp3299 & tmp3300;
    assign tmp3302 = ~tmp57;
    assign tmp3303 = tmp3301 & tmp3302;
    assign tmp3304 = ~tmp1034;
    assign tmp3305 = tmp3303 & tmp3304;
    assign tmp3306 = tmp3305 & tmp2071;
    assign tmp3307 = ~tmp2583;
    assign tmp3308 = tmp3306 & tmp3307;
    assign tmp3309 = tmp3308 & tmp23;
    assign tmp3310 = ~tmp2627;
    assign tmp3311 = tmp3309 & tmp3310;
    assign tmp3312 = tmp3311 & tmp2798;
    assign tmp3313 = ~tmp24;
    assign tmp3314 = tmp3312 & tmp3313;
    assign tmp3315 = {tmp25[255]};
    assign tmp3316 = {tmp29[255]};
    assign tmp3317 = tmp29 - tmp25;
    assign tmp3318 = {tmp3317[256]};
    assign tmp3319 = {tmp25[255]};
    assign tmp3320 = ~tmp3319;
    assign tmp3321 = tmp3318 ^ tmp3320;
    assign tmp3322 = {tmp29[255]};
    assign tmp3323 = ~tmp3322;
    assign tmp3324 = tmp3321 ^ tmp3323;
    assign tmp3325 = tmp25 == tmp29;
    assign tmp3326 = tmp3324 | tmp3325;
    assign tmp3327 = {tmp26[255]};
    assign tmp3328 = {tmp30[255]};
    assign tmp3329 = tmp30 - tmp26;
    assign tmp3330 = {tmp3329[256]};
    assign tmp3331 = {tmp26[255]};
    assign tmp3332 = ~tmp3331;
    assign tmp3333 = tmp3330 ^ tmp3332;
    assign tmp3334 = {tmp30[255]};
    assign tmp3335 = ~tmp3334;
    assign tmp3336 = tmp3333 ^ tmp3335;
    assign tmp3337 = tmp26 == tmp30;
    assign tmp3338 = tmp3336 | tmp3337;
    assign tmp3339 = tmp3326 & tmp3338;
    assign tmp3340 = {tmp27[255]};
    assign tmp3341 = {tmp31[255]};
    assign tmp3342 = tmp31 - tmp27;
    assign tmp3343 = {tmp3342[256]};
    assign tmp3344 = {tmp27[255]};
    assign tmp3345 = ~tmp3344;
    assign tmp3346 = tmp3343 ^ tmp3345;
    assign tmp3347 = {tmp31[255]};
    assign tmp3348 = ~tmp3347;
    assign tmp3349 = tmp3346 ^ tmp3348;
    assign tmp3350 = tmp27 == tmp31;
    assign tmp3351 = tmp3349 | tmp3350;
    assign tmp3352 = tmp3339 & tmp3351;
    assign tmp3353 = {tmp28[255]};
    assign tmp3354 = {tmp32[255]};
    assign tmp3355 = tmp32 - tmp28;
    assign tmp3356 = {tmp3355[256]};
    assign tmp3357 = {tmp28[255]};
    assign tmp3358 = ~tmp3357;
    assign tmp3359 = tmp3356 ^ tmp3358;
    assign tmp3360 = {tmp32[255]};
    assign tmp3361 = ~tmp3360;
    assign tmp3362 = tmp3359 ^ tmp3361;
    assign tmp3363 = tmp28 == tmp32;
    assign tmp3364 = tmp3362 | tmp3363;
    assign tmp3365 = tmp3352 & tmp3364;
    assign tmp3366 = {tmp25[255], tmp25[254], tmp25[253], tmp25[252], tmp25[251], tmp25[250], tmp25[249], tmp25[248], tmp25[247], tmp25[246], tmp25[245], tmp25[244], tmp25[243], tmp25[242], tmp25[241], tmp25[240], tmp25[239], tmp25[238], tmp25[237], tmp25[236], tmp25[235], tmp25[234], tmp25[233], tmp25[232], tmp25[231], tmp25[230], tmp25[229], tmp25[228], tmp25[227], tmp25[226], tmp25[225], tmp25[224], tmp25[223], tmp25[222], tmp25[221], tmp25[220], tmp25[219], tmp25[218], tmp25[217], tmp25[216], tmp25[215], tmp25[214], tmp25[213], tmp25[212], tmp25[211], tmp25[210], tmp25[209], tmp25[208], tmp25[207], tmp25[206], tmp25[205], tmp25[204], tmp25[203], tmp25[202], tmp25[201], tmp25[200], tmp25[199], tmp25[198], tmp25[197], tmp25[196], tmp25[195], tmp25[194], tmp25[193], tmp25[192], tmp25[191], tmp25[190], tmp25[189], tmp25[188], tmp25[187], tmp25[186], tmp25[185], tmp25[184], tmp25[183], tmp25[182], tmp25[181], tmp25[180], tmp25[179], tmp25[178], tmp25[177], tmp25[176], tmp25[175], tmp25[174], tmp25[173], tmp25[172], tmp25[171], tmp25[170], tmp25[169], tmp25[168], tmp25[167], tmp25[166], tmp25[165], tmp25[164], tmp25[163], tmp25[162], tmp25[161], tmp25[160], tmp25[159], tmp25[158], tmp25[157], tmp25[156], tmp25[155], tmp25[154], tmp25[153], tmp25[152], tmp25[151], tmp25[150], tmp25[149], tmp25[148], tmp25[147], tmp25[146], tmp25[145], tmp25[144], tmp25[143], tmp25[142], tmp25[141], tmp25[140], tmp25[139], tmp25[138], tmp25[137], tmp25[136], tmp25[135], tmp25[134], tmp25[133], tmp25[132], tmp25[131], tmp25[130], tmp25[129], tmp25[128], tmp25[127], tmp25[126], tmp25[125], tmp25[124], tmp25[123], tmp25[122], tmp25[121], tmp25[120], tmp25[119], tmp25[118], tmp25[117], tmp25[116], tmp25[115], tmp25[114], tmp25[113], tmp25[112], tmp25[111], tmp25[110], tmp25[109], tmp25[108], tmp25[107], tmp25[106], tmp25[105], tmp25[104], tmp25[103], tmp25[102], tmp25[101], tmp25[100], tmp25[99], tmp25[98], tmp25[97], tmp25[96], tmp25[95], tmp25[94], tmp25[93], tmp25[92], tmp25[91], tmp25[90], tmp25[89], tmp25[88], tmp25[87], tmp25[86], tmp25[85], tmp25[84], tmp25[83], tmp25[82], tmp25[81], tmp25[80], tmp25[79], tmp25[78], tmp25[77], tmp25[76], tmp25[75], tmp25[74], tmp25[73], tmp25[72], tmp25[71], tmp25[70], tmp25[69], tmp25[68], tmp25[67], tmp25[66], tmp25[65], tmp25[64], tmp25[63], tmp25[62], tmp25[61], tmp25[60], tmp25[59], tmp25[58], tmp25[57], tmp25[56], tmp25[55], tmp25[54], tmp25[53], tmp25[52], tmp25[51], tmp25[50], tmp25[49], tmp25[48], tmp25[47], tmp25[46], tmp25[45], tmp25[44], tmp25[43], tmp25[42], tmp25[41], tmp25[40], tmp25[39], tmp25[38], tmp25[37], tmp25[36], tmp25[35], tmp25[34], tmp25[33], tmp25[32], tmp25[31], tmp25[30], tmp25[29], tmp25[28], tmp25[27], tmp25[26], tmp25[25], tmp25[24], tmp25[23], tmp25[22], tmp25[21], tmp25[20], tmp25[19], tmp25[18], tmp25[17], tmp25[16], tmp25[15], tmp25[14], tmp25[13], tmp25[12], tmp25[11], tmp25[10], tmp25[9], tmp25[8], tmp25[7], tmp25[6], tmp25[5], tmp25[4], tmp25[3], tmp25[2], tmp25[1]};
    assign tmp3367 = {tmp3366[254]};
    assign tmp3368 = {tmp3367};
    assign tmp3369 = {tmp3368, tmp3366};
    assign tmp3370 = {tmp3369[255]};
    assign tmp3371 = {tmp29[255]};
    assign tmp3372 = tmp3369 - tmp29;
    assign tmp3373 = {tmp3372[256]};
    assign tmp3374 = {tmp3369[255]};
    assign tmp3375 = ~tmp3374;
    assign tmp3376 = tmp3373 ^ tmp3375;
    assign tmp3377 = {tmp29[255]};
    assign tmp3378 = ~tmp3377;
    assign tmp3379 = tmp3376 ^ tmp3378;
    assign tmp3380 = tmp3365 & tmp3379;
    assign tmp3381 = {tmp26[255], tmp26[254], tmp26[253], tmp26[252], tmp26[251], tmp26[250], tmp26[249], tmp26[248], tmp26[247], tmp26[246], tmp26[245], tmp26[244], tmp26[243], tmp26[242], tmp26[241], tmp26[240], tmp26[239], tmp26[238], tmp26[237], tmp26[236], tmp26[235], tmp26[234], tmp26[233], tmp26[232], tmp26[231], tmp26[230], tmp26[229], tmp26[228], tmp26[227], tmp26[226], tmp26[225], tmp26[224], tmp26[223], tmp26[222], tmp26[221], tmp26[220], tmp26[219], tmp26[218], tmp26[217], tmp26[216], tmp26[215], tmp26[214], tmp26[213], tmp26[212], tmp26[211], tmp26[210], tmp26[209], tmp26[208], tmp26[207], tmp26[206], tmp26[205], tmp26[204], tmp26[203], tmp26[202], tmp26[201], tmp26[200], tmp26[199], tmp26[198], tmp26[197], tmp26[196], tmp26[195], tmp26[194], tmp26[193], tmp26[192], tmp26[191], tmp26[190], tmp26[189], tmp26[188], tmp26[187], tmp26[186], tmp26[185], tmp26[184], tmp26[183], tmp26[182], tmp26[181], tmp26[180], tmp26[179], tmp26[178], tmp26[177], tmp26[176], tmp26[175], tmp26[174], tmp26[173], tmp26[172], tmp26[171], tmp26[170], tmp26[169], tmp26[168], tmp26[167], tmp26[166], tmp26[165], tmp26[164], tmp26[163], tmp26[162], tmp26[161], tmp26[160], tmp26[159], tmp26[158], tmp26[157], tmp26[156], tmp26[155], tmp26[154], tmp26[153], tmp26[152], tmp26[151], tmp26[150], tmp26[149], tmp26[148], tmp26[147], tmp26[146], tmp26[145], tmp26[144], tmp26[143], tmp26[142], tmp26[141], tmp26[140], tmp26[139], tmp26[138], tmp26[137], tmp26[136], tmp26[135], tmp26[134], tmp26[133], tmp26[132], tmp26[131], tmp26[130], tmp26[129], tmp26[128], tmp26[127], tmp26[126], tmp26[125], tmp26[124], tmp26[123], tmp26[122], tmp26[121], tmp26[120], tmp26[119], tmp26[118], tmp26[117], tmp26[116], tmp26[115], tmp26[114], tmp26[113], tmp26[112], tmp26[111], tmp26[110], tmp26[109], tmp26[108], tmp26[107], tmp26[106], tmp26[105], tmp26[104], tmp26[103], tmp26[102], tmp26[101], tmp26[100], tmp26[99], tmp26[98], tmp26[97], tmp26[96], tmp26[95], tmp26[94], tmp26[93], tmp26[92], tmp26[91], tmp26[90], tmp26[89], tmp26[88], tmp26[87], tmp26[86], tmp26[85], tmp26[84], tmp26[83], tmp26[82], tmp26[81], tmp26[80], tmp26[79], tmp26[78], tmp26[77], tmp26[76], tmp26[75], tmp26[74], tmp26[73], tmp26[72], tmp26[71], tmp26[70], tmp26[69], tmp26[68], tmp26[67], tmp26[66], tmp26[65], tmp26[64], tmp26[63], tmp26[62], tmp26[61], tmp26[60], tmp26[59], tmp26[58], tmp26[57], tmp26[56], tmp26[55], tmp26[54], tmp26[53], tmp26[52], tmp26[51], tmp26[50], tmp26[49], tmp26[48], tmp26[47], tmp26[46], tmp26[45], tmp26[44], tmp26[43], tmp26[42], tmp26[41], tmp26[40], tmp26[39], tmp26[38], tmp26[37], tmp26[36], tmp26[35], tmp26[34], tmp26[33], tmp26[32], tmp26[31], tmp26[30], tmp26[29], tmp26[28], tmp26[27], tmp26[26], tmp26[25], tmp26[24], tmp26[23], tmp26[22], tmp26[21], tmp26[20], tmp26[19], tmp26[18], tmp26[17], tmp26[16], tmp26[15], tmp26[14], tmp26[13], tmp26[12], tmp26[11], tmp26[10], tmp26[9], tmp26[8], tmp26[7], tmp26[6], tmp26[5], tmp26[4], tmp26[3], tmp26[2], tmp26[1]};
    assign tmp3382 = {tmp3381[254]};
    assign tmp3383 = {tmp3382};
    assign tmp3384 = {tmp3383, tmp3381};
    assign tmp3385 = {tmp3384[255]};
    assign tmp3386 = {tmp30[255]};
    assign tmp3387 = tmp3384 - tmp30;
    assign tmp3388 = {tmp3387[256]};
    assign tmp3389 = {tmp3384[255]};
    assign tmp3390 = ~tmp3389;
    assign tmp3391 = tmp3388 ^ tmp3390;
    assign tmp3392 = {tmp30[255]};
    assign tmp3393 = ~tmp3392;
    assign tmp3394 = tmp3391 ^ tmp3393;
    assign tmp3395 = tmp3380 & tmp3394;
    assign tmp3396 = {tmp27[255], tmp27[254], tmp27[253], tmp27[252], tmp27[251], tmp27[250], tmp27[249], tmp27[248], tmp27[247], tmp27[246], tmp27[245], tmp27[244], tmp27[243], tmp27[242], tmp27[241], tmp27[240], tmp27[239], tmp27[238], tmp27[237], tmp27[236], tmp27[235], tmp27[234], tmp27[233], tmp27[232], tmp27[231], tmp27[230], tmp27[229], tmp27[228], tmp27[227], tmp27[226], tmp27[225], tmp27[224], tmp27[223], tmp27[222], tmp27[221], tmp27[220], tmp27[219], tmp27[218], tmp27[217], tmp27[216], tmp27[215], tmp27[214], tmp27[213], tmp27[212], tmp27[211], tmp27[210], tmp27[209], tmp27[208], tmp27[207], tmp27[206], tmp27[205], tmp27[204], tmp27[203], tmp27[202], tmp27[201], tmp27[200], tmp27[199], tmp27[198], tmp27[197], tmp27[196], tmp27[195], tmp27[194], tmp27[193], tmp27[192], tmp27[191], tmp27[190], tmp27[189], tmp27[188], tmp27[187], tmp27[186], tmp27[185], tmp27[184], tmp27[183], tmp27[182], tmp27[181], tmp27[180], tmp27[179], tmp27[178], tmp27[177], tmp27[176], tmp27[175], tmp27[174], tmp27[173], tmp27[172], tmp27[171], tmp27[170], tmp27[169], tmp27[168], tmp27[167], tmp27[166], tmp27[165], tmp27[164], tmp27[163], tmp27[162], tmp27[161], tmp27[160], tmp27[159], tmp27[158], tmp27[157], tmp27[156], tmp27[155], tmp27[154], tmp27[153], tmp27[152], tmp27[151], tmp27[150], tmp27[149], tmp27[148], tmp27[147], tmp27[146], tmp27[145], tmp27[144], tmp27[143], tmp27[142], tmp27[141], tmp27[140], tmp27[139], tmp27[138], tmp27[137], tmp27[136], tmp27[135], tmp27[134], tmp27[133], tmp27[132], tmp27[131], tmp27[130], tmp27[129], tmp27[128], tmp27[127], tmp27[126], tmp27[125], tmp27[124], tmp27[123], tmp27[122], tmp27[121], tmp27[120], tmp27[119], tmp27[118], tmp27[117], tmp27[116], tmp27[115], tmp27[114], tmp27[113], tmp27[112], tmp27[111], tmp27[110], tmp27[109], tmp27[108], tmp27[107], tmp27[106], tmp27[105], tmp27[104], tmp27[103], tmp27[102], tmp27[101], tmp27[100], tmp27[99], tmp27[98], tmp27[97], tmp27[96], tmp27[95], tmp27[94], tmp27[93], tmp27[92], tmp27[91], tmp27[90], tmp27[89], tmp27[88], tmp27[87], tmp27[86], tmp27[85], tmp27[84], tmp27[83], tmp27[82], tmp27[81], tmp27[80], tmp27[79], tmp27[78], tmp27[77], tmp27[76], tmp27[75], tmp27[74], tmp27[73], tmp27[72], tmp27[71], tmp27[70], tmp27[69], tmp27[68], tmp27[67], tmp27[66], tmp27[65], tmp27[64], tmp27[63], tmp27[62], tmp27[61], tmp27[60], tmp27[59], tmp27[58], tmp27[57], tmp27[56], tmp27[55], tmp27[54], tmp27[53], tmp27[52], tmp27[51], tmp27[50], tmp27[49], tmp27[48], tmp27[47], tmp27[46], tmp27[45], tmp27[44], tmp27[43], tmp27[42], tmp27[41], tmp27[40], tmp27[39], tmp27[38], tmp27[37], tmp27[36], tmp27[35], tmp27[34], tmp27[33], tmp27[32], tmp27[31], tmp27[30], tmp27[29], tmp27[28], tmp27[27], tmp27[26], tmp27[25], tmp27[24], tmp27[23], tmp27[22], tmp27[21], tmp27[20], tmp27[19], tmp27[18], tmp27[17], tmp27[16], tmp27[15], tmp27[14], tmp27[13], tmp27[12], tmp27[11], tmp27[10], tmp27[9], tmp27[8], tmp27[7], tmp27[6], tmp27[5], tmp27[4], tmp27[3], tmp27[2], tmp27[1]};
    assign tmp3397 = {tmp3396[254]};
    assign tmp3398 = {tmp3397};
    assign tmp3399 = {tmp3398, tmp3396};
    assign tmp3400 = {tmp3399[255]};
    assign tmp3401 = {tmp31[255]};
    assign tmp3402 = tmp3399 - tmp31;
    assign tmp3403 = {tmp3402[256]};
    assign tmp3404 = {tmp3399[255]};
    assign tmp3405 = ~tmp3404;
    assign tmp3406 = tmp3403 ^ tmp3405;
    assign tmp3407 = {tmp31[255]};
    assign tmp3408 = ~tmp3407;
    assign tmp3409 = tmp3406 ^ tmp3408;
    assign tmp3410 = tmp3395 & tmp3409;
    assign tmp3411 = {tmp28[255], tmp28[254], tmp28[253], tmp28[252], tmp28[251], tmp28[250], tmp28[249], tmp28[248], tmp28[247], tmp28[246], tmp28[245], tmp28[244], tmp28[243], tmp28[242], tmp28[241], tmp28[240], tmp28[239], tmp28[238], tmp28[237], tmp28[236], tmp28[235], tmp28[234], tmp28[233], tmp28[232], tmp28[231], tmp28[230], tmp28[229], tmp28[228], tmp28[227], tmp28[226], tmp28[225], tmp28[224], tmp28[223], tmp28[222], tmp28[221], tmp28[220], tmp28[219], tmp28[218], tmp28[217], tmp28[216], tmp28[215], tmp28[214], tmp28[213], tmp28[212], tmp28[211], tmp28[210], tmp28[209], tmp28[208], tmp28[207], tmp28[206], tmp28[205], tmp28[204], tmp28[203], tmp28[202], tmp28[201], tmp28[200], tmp28[199], tmp28[198], tmp28[197], tmp28[196], tmp28[195], tmp28[194], tmp28[193], tmp28[192], tmp28[191], tmp28[190], tmp28[189], tmp28[188], tmp28[187], tmp28[186], tmp28[185], tmp28[184], tmp28[183], tmp28[182], tmp28[181], tmp28[180], tmp28[179], tmp28[178], tmp28[177], tmp28[176], tmp28[175], tmp28[174], tmp28[173], tmp28[172], tmp28[171], tmp28[170], tmp28[169], tmp28[168], tmp28[167], tmp28[166], tmp28[165], tmp28[164], tmp28[163], tmp28[162], tmp28[161], tmp28[160], tmp28[159], tmp28[158], tmp28[157], tmp28[156], tmp28[155], tmp28[154], tmp28[153], tmp28[152], tmp28[151], tmp28[150], tmp28[149], tmp28[148], tmp28[147], tmp28[146], tmp28[145], tmp28[144], tmp28[143], tmp28[142], tmp28[141], tmp28[140], tmp28[139], tmp28[138], tmp28[137], tmp28[136], tmp28[135], tmp28[134], tmp28[133], tmp28[132], tmp28[131], tmp28[130], tmp28[129], tmp28[128], tmp28[127], tmp28[126], tmp28[125], tmp28[124], tmp28[123], tmp28[122], tmp28[121], tmp28[120], tmp28[119], tmp28[118], tmp28[117], tmp28[116], tmp28[115], tmp28[114], tmp28[113], tmp28[112], tmp28[111], tmp28[110], tmp28[109], tmp28[108], tmp28[107], tmp28[106], tmp28[105], tmp28[104], tmp28[103], tmp28[102], tmp28[101], tmp28[100], tmp28[99], tmp28[98], tmp28[97], tmp28[96], tmp28[95], tmp28[94], tmp28[93], tmp28[92], tmp28[91], tmp28[90], tmp28[89], tmp28[88], tmp28[87], tmp28[86], tmp28[85], tmp28[84], tmp28[83], tmp28[82], tmp28[81], tmp28[80], tmp28[79], tmp28[78], tmp28[77], tmp28[76], tmp28[75], tmp28[74], tmp28[73], tmp28[72], tmp28[71], tmp28[70], tmp28[69], tmp28[68], tmp28[67], tmp28[66], tmp28[65], tmp28[64], tmp28[63], tmp28[62], tmp28[61], tmp28[60], tmp28[59], tmp28[58], tmp28[57], tmp28[56], tmp28[55], tmp28[54], tmp28[53], tmp28[52], tmp28[51], tmp28[50], tmp28[49], tmp28[48], tmp28[47], tmp28[46], tmp28[45], tmp28[44], tmp28[43], tmp28[42], tmp28[41], tmp28[40], tmp28[39], tmp28[38], tmp28[37], tmp28[36], tmp28[35], tmp28[34], tmp28[33], tmp28[32], tmp28[31], tmp28[30], tmp28[29], tmp28[28], tmp28[27], tmp28[26], tmp28[25], tmp28[24], tmp28[23], tmp28[22], tmp28[21], tmp28[20], tmp28[19], tmp28[18], tmp28[17], tmp28[16], tmp28[15], tmp28[14], tmp28[13], tmp28[12], tmp28[11], tmp28[10], tmp28[9], tmp28[8], tmp28[7], tmp28[6], tmp28[5], tmp28[4], tmp28[3], tmp28[2], tmp28[1]};
    assign tmp3412 = {tmp3411[254]};
    assign tmp3413 = {tmp3412};
    assign tmp3414 = {tmp3413, tmp3411};
    assign tmp3415 = {tmp3414[255]};
    assign tmp3416 = {tmp32[255]};
    assign tmp3417 = tmp3414 - tmp32;
    assign tmp3418 = {tmp3417[256]};
    assign tmp3419 = {tmp3414[255]};
    assign tmp3420 = ~tmp3419;
    assign tmp3421 = tmp3418 ^ tmp3420;
    assign tmp3422 = {tmp32[255]};
    assign tmp3423 = ~tmp3422;
    assign tmp3424 = tmp3421 ^ tmp3423;
    assign tmp3425 = tmp3410 & tmp3424;
    assign tmp3426 = ~tmp35;
    assign tmp3427 = ~tmp36;
    assign tmp3428 = tmp3426 & tmp3427;
    assign tmp3429 = ~tmp57;
    assign tmp3430 = tmp3428 & tmp3429;
    assign tmp3431 = ~tmp1034;
    assign tmp3432 = tmp3430 & tmp3431;
    assign tmp3433 = tmp3432 & tmp2071;
    assign tmp3434 = ~tmp2583;
    assign tmp3435 = tmp3433 & tmp3434;
    assign tmp3436 = tmp3435 & tmp23;
    assign tmp3437 = ~tmp2627;
    assign tmp3438 = tmp3436 & tmp3437;
    assign tmp3439 = ~tmp2798;
    assign tmp3440 = tmp3438 & tmp3439;
    assign tmp3441 = tmp3440 & tmp3425;
    assign tmp3442 = ~tmp35;
    assign tmp3443 = ~tmp36;
    assign tmp3444 = tmp3442 & tmp3443;
    assign tmp3445 = ~tmp57;
    assign tmp3446 = tmp3444 & tmp3445;
    assign tmp3447 = ~tmp1034;
    assign tmp3448 = tmp3446 & tmp3447;
    assign tmp3449 = tmp3448 & tmp2071;
    assign tmp3450 = ~tmp2583;
    assign tmp3451 = tmp3449 & tmp3450;
    assign tmp3452 = tmp3451 & tmp23;
    assign tmp3453 = ~tmp2627;
    assign tmp3454 = tmp3452 & tmp3453;
    assign tmp3455 = ~tmp2798;
    assign tmp3456 = tmp3454 & tmp3455;
    assign tmp3457 = tmp3456 & tmp3425;
    assign tmp3458 = ~tmp35;
    assign tmp3459 = ~tmp36;
    assign tmp3460 = tmp3458 & tmp3459;
    assign tmp3461 = ~tmp57;
    assign tmp3462 = tmp3460 & tmp3461;
    assign tmp3463 = ~tmp1034;
    assign tmp3464 = tmp3462 & tmp3463;
    assign tmp3465 = tmp3464 & tmp2071;
    assign tmp3466 = ~tmp2583;
    assign tmp3467 = tmp3465 & tmp3466;
    assign tmp3468 = tmp3467 & tmp23;
    assign tmp3469 = ~tmp2627;
    assign tmp3470 = tmp3468 & tmp3469;
    assign tmp3471 = ~tmp2798;
    assign tmp3472 = tmp3470 & tmp3471;
    assign tmp3473 = tmp3472 & tmp3425;
    assign tmp3474 = _ver_out_tmp_16 == tmp29;
    assign tmp3475 = {const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0, const_351_0};
    assign tmp3476 = {tmp3475, const_350_0};
    assign tmp3477 = tmp3476 - tmp29;
    assign tmp3478 = {const_353_0, const_353_0};
    assign tmp3479 = {tmp3478, const_352_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp3480 = tmp3474 ? tmp3479 : tmp3477;
    assign tmp3481 = {tmp25[255]};
    assign tmp3482 = {tmp3481, tmp3481};
    assign tmp3483 = {tmp3482, tmp25};
    assign tmp3484 = {tmp3480[256]};
    assign tmp3485 = {tmp3484};
    assign tmp3486 = {tmp3485, tmp3480};
    assign tmp3487 = tmp3483 + tmp3486;
    assign tmp3488 = {tmp3487[257], tmp3487[256], tmp3487[255], tmp3487[254], tmp3487[253], tmp3487[252], tmp3487[251], tmp3487[250], tmp3487[249], tmp3487[248], tmp3487[247], tmp3487[246], tmp3487[245], tmp3487[244], tmp3487[243], tmp3487[242], tmp3487[241], tmp3487[240], tmp3487[239], tmp3487[238], tmp3487[237], tmp3487[236], tmp3487[235], tmp3487[234], tmp3487[233], tmp3487[232], tmp3487[231], tmp3487[230], tmp3487[229], tmp3487[228], tmp3487[227], tmp3487[226], tmp3487[225], tmp3487[224], tmp3487[223], tmp3487[222], tmp3487[221], tmp3487[220], tmp3487[219], tmp3487[218], tmp3487[217], tmp3487[216], tmp3487[215], tmp3487[214], tmp3487[213], tmp3487[212], tmp3487[211], tmp3487[210], tmp3487[209], tmp3487[208], tmp3487[207], tmp3487[206], tmp3487[205], tmp3487[204], tmp3487[203], tmp3487[202], tmp3487[201], tmp3487[200], tmp3487[199], tmp3487[198], tmp3487[197], tmp3487[196], tmp3487[195], tmp3487[194], tmp3487[193], tmp3487[192], tmp3487[191], tmp3487[190], tmp3487[189], tmp3487[188], tmp3487[187], tmp3487[186], tmp3487[185], tmp3487[184], tmp3487[183], tmp3487[182], tmp3487[181], tmp3487[180], tmp3487[179], tmp3487[178], tmp3487[177], tmp3487[176], tmp3487[175], tmp3487[174], tmp3487[173], tmp3487[172], tmp3487[171], tmp3487[170], tmp3487[169], tmp3487[168], tmp3487[167], tmp3487[166], tmp3487[165], tmp3487[164], tmp3487[163], tmp3487[162], tmp3487[161], tmp3487[160], tmp3487[159], tmp3487[158], tmp3487[157], tmp3487[156], tmp3487[155], tmp3487[154], tmp3487[153], tmp3487[152], tmp3487[151], tmp3487[150], tmp3487[149], tmp3487[148], tmp3487[147], tmp3487[146], tmp3487[145], tmp3487[144], tmp3487[143], tmp3487[142], tmp3487[141], tmp3487[140], tmp3487[139], tmp3487[138], tmp3487[137], tmp3487[136], tmp3487[135], tmp3487[134], tmp3487[133], tmp3487[132], tmp3487[131], tmp3487[130], tmp3487[129], tmp3487[128], tmp3487[127], tmp3487[126], tmp3487[125], tmp3487[124], tmp3487[123], tmp3487[122], tmp3487[121], tmp3487[120], tmp3487[119], tmp3487[118], tmp3487[117], tmp3487[116], tmp3487[115], tmp3487[114], tmp3487[113], tmp3487[112], tmp3487[111], tmp3487[110], tmp3487[109], tmp3487[108], tmp3487[107], tmp3487[106], tmp3487[105], tmp3487[104], tmp3487[103], tmp3487[102], tmp3487[101], tmp3487[100], tmp3487[99], tmp3487[98], tmp3487[97], tmp3487[96], tmp3487[95], tmp3487[94], tmp3487[93], tmp3487[92], tmp3487[91], tmp3487[90], tmp3487[89], tmp3487[88], tmp3487[87], tmp3487[86], tmp3487[85], tmp3487[84], tmp3487[83], tmp3487[82], tmp3487[81], tmp3487[80], tmp3487[79], tmp3487[78], tmp3487[77], tmp3487[76], tmp3487[75], tmp3487[74], tmp3487[73], tmp3487[72], tmp3487[71], tmp3487[70], tmp3487[69], tmp3487[68], tmp3487[67], tmp3487[66], tmp3487[65], tmp3487[64], tmp3487[63], tmp3487[62], tmp3487[61], tmp3487[60], tmp3487[59], tmp3487[58], tmp3487[57], tmp3487[56], tmp3487[55], tmp3487[54], tmp3487[53], tmp3487[52], tmp3487[51], tmp3487[50], tmp3487[49], tmp3487[48], tmp3487[47], tmp3487[46], tmp3487[45], tmp3487[44], tmp3487[43], tmp3487[42], tmp3487[41], tmp3487[40], tmp3487[39], tmp3487[38], tmp3487[37], tmp3487[36], tmp3487[35], tmp3487[34], tmp3487[33], tmp3487[32], tmp3487[31], tmp3487[30], tmp3487[29], tmp3487[28], tmp3487[27], tmp3487[26], tmp3487[25], tmp3487[24], tmp3487[23], tmp3487[22], tmp3487[21], tmp3487[20], tmp3487[19], tmp3487[18], tmp3487[17], tmp3487[16], tmp3487[15], tmp3487[14], tmp3487[13], tmp3487[12], tmp3487[11], tmp3487[10], tmp3487[9], tmp3487[8], tmp3487[7], tmp3487[6], tmp3487[5], tmp3487[4], tmp3487[3], tmp3487[2], tmp3487[1], tmp3487[0]};
    assign tmp3489 = {tmp3488[255], tmp3488[254], tmp3488[253], tmp3488[252], tmp3488[251], tmp3488[250], tmp3488[249], tmp3488[248], tmp3488[247], tmp3488[246], tmp3488[245], tmp3488[244], tmp3488[243], tmp3488[242], tmp3488[241], tmp3488[240], tmp3488[239], tmp3488[238], tmp3488[237], tmp3488[236], tmp3488[235], tmp3488[234], tmp3488[233], tmp3488[232], tmp3488[231], tmp3488[230], tmp3488[229], tmp3488[228], tmp3488[227], tmp3488[226], tmp3488[225], tmp3488[224], tmp3488[223], tmp3488[222], tmp3488[221], tmp3488[220], tmp3488[219], tmp3488[218], tmp3488[217], tmp3488[216], tmp3488[215], tmp3488[214], tmp3488[213], tmp3488[212], tmp3488[211], tmp3488[210], tmp3488[209], tmp3488[208], tmp3488[207], tmp3488[206], tmp3488[205], tmp3488[204], tmp3488[203], tmp3488[202], tmp3488[201], tmp3488[200], tmp3488[199], tmp3488[198], tmp3488[197], tmp3488[196], tmp3488[195], tmp3488[194], tmp3488[193], tmp3488[192], tmp3488[191], tmp3488[190], tmp3488[189], tmp3488[188], tmp3488[187], tmp3488[186], tmp3488[185], tmp3488[184], tmp3488[183], tmp3488[182], tmp3488[181], tmp3488[180], tmp3488[179], tmp3488[178], tmp3488[177], tmp3488[176], tmp3488[175], tmp3488[174], tmp3488[173], tmp3488[172], tmp3488[171], tmp3488[170], tmp3488[169], tmp3488[168], tmp3488[167], tmp3488[166], tmp3488[165], tmp3488[164], tmp3488[163], tmp3488[162], tmp3488[161], tmp3488[160], tmp3488[159], tmp3488[158], tmp3488[157], tmp3488[156], tmp3488[155], tmp3488[154], tmp3488[153], tmp3488[152], tmp3488[151], tmp3488[150], tmp3488[149], tmp3488[148], tmp3488[147], tmp3488[146], tmp3488[145], tmp3488[144], tmp3488[143], tmp3488[142], tmp3488[141], tmp3488[140], tmp3488[139], tmp3488[138], tmp3488[137], tmp3488[136], tmp3488[135], tmp3488[134], tmp3488[133], tmp3488[132], tmp3488[131], tmp3488[130], tmp3488[129], tmp3488[128], tmp3488[127], tmp3488[126], tmp3488[125], tmp3488[124], tmp3488[123], tmp3488[122], tmp3488[121], tmp3488[120], tmp3488[119], tmp3488[118], tmp3488[117], tmp3488[116], tmp3488[115], tmp3488[114], tmp3488[113], tmp3488[112], tmp3488[111], tmp3488[110], tmp3488[109], tmp3488[108], tmp3488[107], tmp3488[106], tmp3488[105], tmp3488[104], tmp3488[103], tmp3488[102], tmp3488[101], tmp3488[100], tmp3488[99], tmp3488[98], tmp3488[97], tmp3488[96], tmp3488[95], tmp3488[94], tmp3488[93], tmp3488[92], tmp3488[91], tmp3488[90], tmp3488[89], tmp3488[88], tmp3488[87], tmp3488[86], tmp3488[85], tmp3488[84], tmp3488[83], tmp3488[82], tmp3488[81], tmp3488[80], tmp3488[79], tmp3488[78], tmp3488[77], tmp3488[76], tmp3488[75], tmp3488[74], tmp3488[73], tmp3488[72], tmp3488[71], tmp3488[70], tmp3488[69], tmp3488[68], tmp3488[67], tmp3488[66], tmp3488[65], tmp3488[64], tmp3488[63], tmp3488[62], tmp3488[61], tmp3488[60], tmp3488[59], tmp3488[58], tmp3488[57], tmp3488[56], tmp3488[55], tmp3488[54], tmp3488[53], tmp3488[52], tmp3488[51], tmp3488[50], tmp3488[49], tmp3488[48], tmp3488[47], tmp3488[46], tmp3488[45], tmp3488[44], tmp3488[43], tmp3488[42], tmp3488[41], tmp3488[40], tmp3488[39], tmp3488[38], tmp3488[37], tmp3488[36], tmp3488[35], tmp3488[34], tmp3488[33], tmp3488[32], tmp3488[31], tmp3488[30], tmp3488[29], tmp3488[28], tmp3488[27], tmp3488[26], tmp3488[25], tmp3488[24], tmp3488[23], tmp3488[22], tmp3488[21], tmp3488[20], tmp3488[19], tmp3488[18], tmp3488[17], tmp3488[16], tmp3488[15], tmp3488[14], tmp3488[13], tmp3488[12], tmp3488[11], tmp3488[10], tmp3488[9], tmp3488[8], tmp3488[7], tmp3488[6], tmp3488[5], tmp3488[4], tmp3488[3], tmp3488[2], tmp3488[1], tmp3488[0]};
    assign tmp3490 = {const_354_0};
    assign tmp3491 = {tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490, tmp3490};
    assign tmp3492 = {tmp3491, const_354_0};
    assign tmp3493 = {tmp25[255]};
    assign tmp3494 = tmp3492 - tmp25;
    assign tmp3495 = {tmp3494[256]};
    assign tmp3496 = {tmp3492[255]};
    assign tmp3497 = ~tmp3496;
    assign tmp3498 = tmp3495 ^ tmp3497;
    assign tmp3499 = {tmp25[255]};
    assign tmp3500 = ~tmp3499;
    assign tmp3501 = tmp3498 ^ tmp3500;
    assign tmp3502 = {const_355_0};
    assign tmp3503 = {tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502, tmp3502};
    assign tmp3504 = {tmp3503, const_355_0};
    assign tmp3505 = {tmp3480[256]};
    assign tmp3506 = tmp3504 - tmp3480;
    assign tmp3507 = {tmp3506[257]};
    assign tmp3508 = {tmp3504[256]};
    assign tmp3509 = ~tmp3508;
    assign tmp3510 = tmp3507 ^ tmp3509;
    assign tmp3511 = {tmp3480[256]};
    assign tmp3512 = ~tmp3511;
    assign tmp3513 = tmp3510 ^ tmp3512;
    assign tmp3514 = tmp3501 & tmp3513;
    assign tmp3515 = {tmp3489[255]};
    assign tmp3516 = {const_356_0};
    assign tmp3517 = {tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516, tmp3516};
    assign tmp3518 = {tmp3517, const_356_0};
    assign tmp3519 = tmp3489 - tmp3518;
    assign tmp3520 = {tmp3519[256]};
    assign tmp3521 = {tmp3489[255]};
    assign tmp3522 = ~tmp3521;
    assign tmp3523 = tmp3520 ^ tmp3522;
    assign tmp3524 = {tmp3518[255]};
    assign tmp3525 = ~tmp3524;
    assign tmp3526 = tmp3523 ^ tmp3525;
    assign tmp3527 = tmp3489 == tmp3518;
    assign tmp3528 = tmp3526 | tmp3527;
    assign tmp3529 = tmp3514 & tmp3528;
    assign tmp3530 = {tmp25[255]};
    assign tmp3531 = {const_357_0};
    assign tmp3532 = {tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531, tmp3531};
    assign tmp3533 = {tmp3532, const_357_0};
    assign tmp3534 = tmp25 - tmp3533;
    assign tmp3535 = {tmp3534[256]};
    assign tmp3536 = {tmp25[255]};
    assign tmp3537 = ~tmp3536;
    assign tmp3538 = tmp3535 ^ tmp3537;
    assign tmp3539 = {tmp3533[255]};
    assign tmp3540 = ~tmp3539;
    assign tmp3541 = tmp3538 ^ tmp3540;
    assign tmp3542 = {tmp3480[256]};
    assign tmp3543 = {const_358_0};
    assign tmp3544 = {tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543, tmp3543};
    assign tmp3545 = {tmp3544, const_358_0};
    assign tmp3546 = tmp3480 - tmp3545;
    assign tmp3547 = {tmp3546[257]};
    assign tmp3548 = {tmp3480[256]};
    assign tmp3549 = ~tmp3548;
    assign tmp3550 = tmp3547 ^ tmp3549;
    assign tmp3551 = {tmp3545[256]};
    assign tmp3552 = ~tmp3551;
    assign tmp3553 = tmp3550 ^ tmp3552;
    assign tmp3554 = tmp3541 & tmp3553;
    assign tmp3555 = {const_359_0};
    assign tmp3556 = {tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555, tmp3555};
    assign tmp3557 = {tmp3556, const_359_0};
    assign tmp3558 = {tmp3489[255]};
    assign tmp3559 = tmp3557 - tmp3489;
    assign tmp3560 = {tmp3559[256]};
    assign tmp3561 = {tmp3557[255]};
    assign tmp3562 = ~tmp3561;
    assign tmp3563 = tmp3560 ^ tmp3562;
    assign tmp3564 = {tmp3489[255]};
    assign tmp3565 = ~tmp3564;
    assign tmp3566 = tmp3563 ^ tmp3565;
    assign tmp3567 = tmp3557 == tmp3489;
    assign tmp3568 = tmp3566 | tmp3567;
    assign tmp3569 = tmp3554 & tmp3568;
    assign tmp3570 = tmp3529 ? const_360_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp3489;
    assign tmp3571 = tmp3569 ? _ver_out_tmp_39 : tmp3570;
    assign tmp3572 = ~tmp35;
    assign tmp3573 = ~tmp36;
    assign tmp3574 = tmp3572 & tmp3573;
    assign tmp3575 = ~tmp57;
    assign tmp3576 = tmp3574 & tmp3575;
    assign tmp3577 = ~tmp1034;
    assign tmp3578 = tmp3576 & tmp3577;
    assign tmp3579 = tmp3578 & tmp2071;
    assign tmp3580 = ~tmp2583;
    assign tmp3581 = tmp3579 & tmp3580;
    assign tmp3582 = tmp3581 & tmp23;
    assign tmp3583 = ~tmp2627;
    assign tmp3584 = tmp3582 & tmp3583;
    assign tmp3585 = ~tmp2798;
    assign tmp3586 = tmp3584 & tmp3585;
    assign tmp3587 = tmp3586 & tmp3425;
    assign tmp3588 = ~tmp35;
    assign tmp3589 = ~tmp36;
    assign tmp3590 = tmp3588 & tmp3589;
    assign tmp3591 = ~tmp57;
    assign tmp3592 = tmp3590 & tmp3591;
    assign tmp3593 = ~tmp1034;
    assign tmp3594 = tmp3592 & tmp3593;
    assign tmp3595 = tmp3594 & tmp2071;
    assign tmp3596 = ~tmp2583;
    assign tmp3597 = tmp3595 & tmp3596;
    assign tmp3598 = tmp3597 & tmp23;
    assign tmp3599 = ~tmp2627;
    assign tmp3600 = tmp3598 & tmp3599;
    assign tmp3601 = ~tmp2798;
    assign tmp3602 = tmp3600 & tmp3601;
    assign tmp3603 = tmp3602 & tmp3425;
    assign tmp3604 = _ver_out_tmp_79 == tmp30;
    assign tmp3605 = {const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0, const_364_0};
    assign tmp3606 = {tmp3605, const_363_0};
    assign tmp3607 = tmp3606 - tmp30;
    assign tmp3608 = {const_366_0, const_366_0};
    assign tmp3609 = {tmp3608, const_365_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp3610 = tmp3604 ? tmp3609 : tmp3607;
    assign tmp3611 = {tmp26[255]};
    assign tmp3612 = {tmp3611, tmp3611};
    assign tmp3613 = {tmp3612, tmp26};
    assign tmp3614 = {tmp3610[256]};
    assign tmp3615 = {tmp3614};
    assign tmp3616 = {tmp3615, tmp3610};
    assign tmp3617 = tmp3613 + tmp3616;
    assign tmp3618 = {tmp3617[257], tmp3617[256], tmp3617[255], tmp3617[254], tmp3617[253], tmp3617[252], tmp3617[251], tmp3617[250], tmp3617[249], tmp3617[248], tmp3617[247], tmp3617[246], tmp3617[245], tmp3617[244], tmp3617[243], tmp3617[242], tmp3617[241], tmp3617[240], tmp3617[239], tmp3617[238], tmp3617[237], tmp3617[236], tmp3617[235], tmp3617[234], tmp3617[233], tmp3617[232], tmp3617[231], tmp3617[230], tmp3617[229], tmp3617[228], tmp3617[227], tmp3617[226], tmp3617[225], tmp3617[224], tmp3617[223], tmp3617[222], tmp3617[221], tmp3617[220], tmp3617[219], tmp3617[218], tmp3617[217], tmp3617[216], tmp3617[215], tmp3617[214], tmp3617[213], tmp3617[212], tmp3617[211], tmp3617[210], tmp3617[209], tmp3617[208], tmp3617[207], tmp3617[206], tmp3617[205], tmp3617[204], tmp3617[203], tmp3617[202], tmp3617[201], tmp3617[200], tmp3617[199], tmp3617[198], tmp3617[197], tmp3617[196], tmp3617[195], tmp3617[194], tmp3617[193], tmp3617[192], tmp3617[191], tmp3617[190], tmp3617[189], tmp3617[188], tmp3617[187], tmp3617[186], tmp3617[185], tmp3617[184], tmp3617[183], tmp3617[182], tmp3617[181], tmp3617[180], tmp3617[179], tmp3617[178], tmp3617[177], tmp3617[176], tmp3617[175], tmp3617[174], tmp3617[173], tmp3617[172], tmp3617[171], tmp3617[170], tmp3617[169], tmp3617[168], tmp3617[167], tmp3617[166], tmp3617[165], tmp3617[164], tmp3617[163], tmp3617[162], tmp3617[161], tmp3617[160], tmp3617[159], tmp3617[158], tmp3617[157], tmp3617[156], tmp3617[155], tmp3617[154], tmp3617[153], tmp3617[152], tmp3617[151], tmp3617[150], tmp3617[149], tmp3617[148], tmp3617[147], tmp3617[146], tmp3617[145], tmp3617[144], tmp3617[143], tmp3617[142], tmp3617[141], tmp3617[140], tmp3617[139], tmp3617[138], tmp3617[137], tmp3617[136], tmp3617[135], tmp3617[134], tmp3617[133], tmp3617[132], tmp3617[131], tmp3617[130], tmp3617[129], tmp3617[128], tmp3617[127], tmp3617[126], tmp3617[125], tmp3617[124], tmp3617[123], tmp3617[122], tmp3617[121], tmp3617[120], tmp3617[119], tmp3617[118], tmp3617[117], tmp3617[116], tmp3617[115], tmp3617[114], tmp3617[113], tmp3617[112], tmp3617[111], tmp3617[110], tmp3617[109], tmp3617[108], tmp3617[107], tmp3617[106], tmp3617[105], tmp3617[104], tmp3617[103], tmp3617[102], tmp3617[101], tmp3617[100], tmp3617[99], tmp3617[98], tmp3617[97], tmp3617[96], tmp3617[95], tmp3617[94], tmp3617[93], tmp3617[92], tmp3617[91], tmp3617[90], tmp3617[89], tmp3617[88], tmp3617[87], tmp3617[86], tmp3617[85], tmp3617[84], tmp3617[83], tmp3617[82], tmp3617[81], tmp3617[80], tmp3617[79], tmp3617[78], tmp3617[77], tmp3617[76], tmp3617[75], tmp3617[74], tmp3617[73], tmp3617[72], tmp3617[71], tmp3617[70], tmp3617[69], tmp3617[68], tmp3617[67], tmp3617[66], tmp3617[65], tmp3617[64], tmp3617[63], tmp3617[62], tmp3617[61], tmp3617[60], tmp3617[59], tmp3617[58], tmp3617[57], tmp3617[56], tmp3617[55], tmp3617[54], tmp3617[53], tmp3617[52], tmp3617[51], tmp3617[50], tmp3617[49], tmp3617[48], tmp3617[47], tmp3617[46], tmp3617[45], tmp3617[44], tmp3617[43], tmp3617[42], tmp3617[41], tmp3617[40], tmp3617[39], tmp3617[38], tmp3617[37], tmp3617[36], tmp3617[35], tmp3617[34], tmp3617[33], tmp3617[32], tmp3617[31], tmp3617[30], tmp3617[29], tmp3617[28], tmp3617[27], tmp3617[26], tmp3617[25], tmp3617[24], tmp3617[23], tmp3617[22], tmp3617[21], tmp3617[20], tmp3617[19], tmp3617[18], tmp3617[17], tmp3617[16], tmp3617[15], tmp3617[14], tmp3617[13], tmp3617[12], tmp3617[11], tmp3617[10], tmp3617[9], tmp3617[8], tmp3617[7], tmp3617[6], tmp3617[5], tmp3617[4], tmp3617[3], tmp3617[2], tmp3617[1], tmp3617[0]};
    assign tmp3619 = {tmp3618[255], tmp3618[254], tmp3618[253], tmp3618[252], tmp3618[251], tmp3618[250], tmp3618[249], tmp3618[248], tmp3618[247], tmp3618[246], tmp3618[245], tmp3618[244], tmp3618[243], tmp3618[242], tmp3618[241], tmp3618[240], tmp3618[239], tmp3618[238], tmp3618[237], tmp3618[236], tmp3618[235], tmp3618[234], tmp3618[233], tmp3618[232], tmp3618[231], tmp3618[230], tmp3618[229], tmp3618[228], tmp3618[227], tmp3618[226], tmp3618[225], tmp3618[224], tmp3618[223], tmp3618[222], tmp3618[221], tmp3618[220], tmp3618[219], tmp3618[218], tmp3618[217], tmp3618[216], tmp3618[215], tmp3618[214], tmp3618[213], tmp3618[212], tmp3618[211], tmp3618[210], tmp3618[209], tmp3618[208], tmp3618[207], tmp3618[206], tmp3618[205], tmp3618[204], tmp3618[203], tmp3618[202], tmp3618[201], tmp3618[200], tmp3618[199], tmp3618[198], tmp3618[197], tmp3618[196], tmp3618[195], tmp3618[194], tmp3618[193], tmp3618[192], tmp3618[191], tmp3618[190], tmp3618[189], tmp3618[188], tmp3618[187], tmp3618[186], tmp3618[185], tmp3618[184], tmp3618[183], tmp3618[182], tmp3618[181], tmp3618[180], tmp3618[179], tmp3618[178], tmp3618[177], tmp3618[176], tmp3618[175], tmp3618[174], tmp3618[173], tmp3618[172], tmp3618[171], tmp3618[170], tmp3618[169], tmp3618[168], tmp3618[167], tmp3618[166], tmp3618[165], tmp3618[164], tmp3618[163], tmp3618[162], tmp3618[161], tmp3618[160], tmp3618[159], tmp3618[158], tmp3618[157], tmp3618[156], tmp3618[155], tmp3618[154], tmp3618[153], tmp3618[152], tmp3618[151], tmp3618[150], tmp3618[149], tmp3618[148], tmp3618[147], tmp3618[146], tmp3618[145], tmp3618[144], tmp3618[143], tmp3618[142], tmp3618[141], tmp3618[140], tmp3618[139], tmp3618[138], tmp3618[137], tmp3618[136], tmp3618[135], tmp3618[134], tmp3618[133], tmp3618[132], tmp3618[131], tmp3618[130], tmp3618[129], tmp3618[128], tmp3618[127], tmp3618[126], tmp3618[125], tmp3618[124], tmp3618[123], tmp3618[122], tmp3618[121], tmp3618[120], tmp3618[119], tmp3618[118], tmp3618[117], tmp3618[116], tmp3618[115], tmp3618[114], tmp3618[113], tmp3618[112], tmp3618[111], tmp3618[110], tmp3618[109], tmp3618[108], tmp3618[107], tmp3618[106], tmp3618[105], tmp3618[104], tmp3618[103], tmp3618[102], tmp3618[101], tmp3618[100], tmp3618[99], tmp3618[98], tmp3618[97], tmp3618[96], tmp3618[95], tmp3618[94], tmp3618[93], tmp3618[92], tmp3618[91], tmp3618[90], tmp3618[89], tmp3618[88], tmp3618[87], tmp3618[86], tmp3618[85], tmp3618[84], tmp3618[83], tmp3618[82], tmp3618[81], tmp3618[80], tmp3618[79], tmp3618[78], tmp3618[77], tmp3618[76], tmp3618[75], tmp3618[74], tmp3618[73], tmp3618[72], tmp3618[71], tmp3618[70], tmp3618[69], tmp3618[68], tmp3618[67], tmp3618[66], tmp3618[65], tmp3618[64], tmp3618[63], tmp3618[62], tmp3618[61], tmp3618[60], tmp3618[59], tmp3618[58], tmp3618[57], tmp3618[56], tmp3618[55], tmp3618[54], tmp3618[53], tmp3618[52], tmp3618[51], tmp3618[50], tmp3618[49], tmp3618[48], tmp3618[47], tmp3618[46], tmp3618[45], tmp3618[44], tmp3618[43], tmp3618[42], tmp3618[41], tmp3618[40], tmp3618[39], tmp3618[38], tmp3618[37], tmp3618[36], tmp3618[35], tmp3618[34], tmp3618[33], tmp3618[32], tmp3618[31], tmp3618[30], tmp3618[29], tmp3618[28], tmp3618[27], tmp3618[26], tmp3618[25], tmp3618[24], tmp3618[23], tmp3618[22], tmp3618[21], tmp3618[20], tmp3618[19], tmp3618[18], tmp3618[17], tmp3618[16], tmp3618[15], tmp3618[14], tmp3618[13], tmp3618[12], tmp3618[11], tmp3618[10], tmp3618[9], tmp3618[8], tmp3618[7], tmp3618[6], tmp3618[5], tmp3618[4], tmp3618[3], tmp3618[2], tmp3618[1], tmp3618[0]};
    assign tmp3620 = {const_367_0};
    assign tmp3621 = {tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620, tmp3620};
    assign tmp3622 = {tmp3621, const_367_0};
    assign tmp3623 = {tmp26[255]};
    assign tmp3624 = tmp3622 - tmp26;
    assign tmp3625 = {tmp3624[256]};
    assign tmp3626 = {tmp3622[255]};
    assign tmp3627 = ~tmp3626;
    assign tmp3628 = tmp3625 ^ tmp3627;
    assign tmp3629 = {tmp26[255]};
    assign tmp3630 = ~tmp3629;
    assign tmp3631 = tmp3628 ^ tmp3630;
    assign tmp3632 = {const_368_0};
    assign tmp3633 = {tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632, tmp3632};
    assign tmp3634 = {tmp3633, const_368_0};
    assign tmp3635 = {tmp3610[256]};
    assign tmp3636 = tmp3634 - tmp3610;
    assign tmp3637 = {tmp3636[257]};
    assign tmp3638 = {tmp3634[256]};
    assign tmp3639 = ~tmp3638;
    assign tmp3640 = tmp3637 ^ tmp3639;
    assign tmp3641 = {tmp3610[256]};
    assign tmp3642 = ~tmp3641;
    assign tmp3643 = tmp3640 ^ tmp3642;
    assign tmp3644 = tmp3631 & tmp3643;
    assign tmp3645 = {tmp3619[255]};
    assign tmp3646 = {const_369_0};
    assign tmp3647 = {tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646, tmp3646};
    assign tmp3648 = {tmp3647, const_369_0};
    assign tmp3649 = tmp3619 - tmp3648;
    assign tmp3650 = {tmp3649[256]};
    assign tmp3651 = {tmp3619[255]};
    assign tmp3652 = ~tmp3651;
    assign tmp3653 = tmp3650 ^ tmp3652;
    assign tmp3654 = {tmp3648[255]};
    assign tmp3655 = ~tmp3654;
    assign tmp3656 = tmp3653 ^ tmp3655;
    assign tmp3657 = tmp3619 == tmp3648;
    assign tmp3658 = tmp3656 | tmp3657;
    assign tmp3659 = tmp3644 & tmp3658;
    assign tmp3660 = {tmp26[255]};
    assign tmp3661 = {const_370_0};
    assign tmp3662 = {tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661, tmp3661};
    assign tmp3663 = {tmp3662, const_370_0};
    assign tmp3664 = tmp26 - tmp3663;
    assign tmp3665 = {tmp3664[256]};
    assign tmp3666 = {tmp26[255]};
    assign tmp3667 = ~tmp3666;
    assign tmp3668 = tmp3665 ^ tmp3667;
    assign tmp3669 = {tmp3663[255]};
    assign tmp3670 = ~tmp3669;
    assign tmp3671 = tmp3668 ^ tmp3670;
    assign tmp3672 = {tmp3610[256]};
    assign tmp3673 = {const_371_0};
    assign tmp3674 = {tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673, tmp3673};
    assign tmp3675 = {tmp3674, const_371_0};
    assign tmp3676 = tmp3610 - tmp3675;
    assign tmp3677 = {tmp3676[257]};
    assign tmp3678 = {tmp3610[256]};
    assign tmp3679 = ~tmp3678;
    assign tmp3680 = tmp3677 ^ tmp3679;
    assign tmp3681 = {tmp3675[256]};
    assign tmp3682 = ~tmp3681;
    assign tmp3683 = tmp3680 ^ tmp3682;
    assign tmp3684 = tmp3671 & tmp3683;
    assign tmp3685 = {const_372_0};
    assign tmp3686 = {tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685, tmp3685};
    assign tmp3687 = {tmp3686, const_372_0};
    assign tmp3688 = {tmp3619[255]};
    assign tmp3689 = tmp3687 - tmp3619;
    assign tmp3690 = {tmp3689[256]};
    assign tmp3691 = {tmp3687[255]};
    assign tmp3692 = ~tmp3691;
    assign tmp3693 = tmp3690 ^ tmp3692;
    assign tmp3694 = {tmp3619[255]};
    assign tmp3695 = ~tmp3694;
    assign tmp3696 = tmp3693 ^ tmp3695;
    assign tmp3697 = tmp3687 == tmp3619;
    assign tmp3698 = tmp3696 | tmp3697;
    assign tmp3699 = tmp3684 & tmp3698;
    assign tmp3700 = tmp3659 ? const_373_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp3619;
    assign tmp3701 = tmp3699 ? _ver_out_tmp_81 : tmp3700;
    assign tmp3702 = ~tmp35;
    assign tmp3703 = ~tmp36;
    assign tmp3704 = tmp3702 & tmp3703;
    assign tmp3705 = ~tmp57;
    assign tmp3706 = tmp3704 & tmp3705;
    assign tmp3707 = ~tmp1034;
    assign tmp3708 = tmp3706 & tmp3707;
    assign tmp3709 = tmp3708 & tmp2071;
    assign tmp3710 = ~tmp2583;
    assign tmp3711 = tmp3709 & tmp3710;
    assign tmp3712 = tmp3711 & tmp23;
    assign tmp3713 = ~tmp2627;
    assign tmp3714 = tmp3712 & tmp3713;
    assign tmp3715 = ~tmp2798;
    assign tmp3716 = tmp3714 & tmp3715;
    assign tmp3717 = tmp3716 & tmp3425;
    assign tmp3718 = ~tmp35;
    assign tmp3719 = ~tmp36;
    assign tmp3720 = tmp3718 & tmp3719;
    assign tmp3721 = ~tmp57;
    assign tmp3722 = tmp3720 & tmp3721;
    assign tmp3723 = ~tmp1034;
    assign tmp3724 = tmp3722 & tmp3723;
    assign tmp3725 = tmp3724 & tmp2071;
    assign tmp3726 = ~tmp2583;
    assign tmp3727 = tmp3725 & tmp3726;
    assign tmp3728 = tmp3727 & tmp23;
    assign tmp3729 = ~tmp2627;
    assign tmp3730 = tmp3728 & tmp3729;
    assign tmp3731 = ~tmp2798;
    assign tmp3732 = tmp3730 & tmp3731;
    assign tmp3733 = tmp3732 & tmp3425;
    assign tmp3734 = _ver_out_tmp_82 == tmp31;
    assign tmp3735 = {const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0, const_377_0};
    assign tmp3736 = {tmp3735, const_376_0};
    assign tmp3737 = tmp3736 - tmp31;
    assign tmp3738 = {const_379_0, const_379_0};
    assign tmp3739 = {tmp3738, const_378_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp3740 = tmp3734 ? tmp3739 : tmp3737;
    assign tmp3741 = {tmp27[255]};
    assign tmp3742 = {tmp3741, tmp3741};
    assign tmp3743 = {tmp3742, tmp27};
    assign tmp3744 = {tmp3740[256]};
    assign tmp3745 = {tmp3744};
    assign tmp3746 = {tmp3745, tmp3740};
    assign tmp3747 = tmp3743 + tmp3746;
    assign tmp3748 = {tmp3747[257], tmp3747[256], tmp3747[255], tmp3747[254], tmp3747[253], tmp3747[252], tmp3747[251], tmp3747[250], tmp3747[249], tmp3747[248], tmp3747[247], tmp3747[246], tmp3747[245], tmp3747[244], tmp3747[243], tmp3747[242], tmp3747[241], tmp3747[240], tmp3747[239], tmp3747[238], tmp3747[237], tmp3747[236], tmp3747[235], tmp3747[234], tmp3747[233], tmp3747[232], tmp3747[231], tmp3747[230], tmp3747[229], tmp3747[228], tmp3747[227], tmp3747[226], tmp3747[225], tmp3747[224], tmp3747[223], tmp3747[222], tmp3747[221], tmp3747[220], tmp3747[219], tmp3747[218], tmp3747[217], tmp3747[216], tmp3747[215], tmp3747[214], tmp3747[213], tmp3747[212], tmp3747[211], tmp3747[210], tmp3747[209], tmp3747[208], tmp3747[207], tmp3747[206], tmp3747[205], tmp3747[204], tmp3747[203], tmp3747[202], tmp3747[201], tmp3747[200], tmp3747[199], tmp3747[198], tmp3747[197], tmp3747[196], tmp3747[195], tmp3747[194], tmp3747[193], tmp3747[192], tmp3747[191], tmp3747[190], tmp3747[189], tmp3747[188], tmp3747[187], tmp3747[186], tmp3747[185], tmp3747[184], tmp3747[183], tmp3747[182], tmp3747[181], tmp3747[180], tmp3747[179], tmp3747[178], tmp3747[177], tmp3747[176], tmp3747[175], tmp3747[174], tmp3747[173], tmp3747[172], tmp3747[171], tmp3747[170], tmp3747[169], tmp3747[168], tmp3747[167], tmp3747[166], tmp3747[165], tmp3747[164], tmp3747[163], tmp3747[162], tmp3747[161], tmp3747[160], tmp3747[159], tmp3747[158], tmp3747[157], tmp3747[156], tmp3747[155], tmp3747[154], tmp3747[153], tmp3747[152], tmp3747[151], tmp3747[150], tmp3747[149], tmp3747[148], tmp3747[147], tmp3747[146], tmp3747[145], tmp3747[144], tmp3747[143], tmp3747[142], tmp3747[141], tmp3747[140], tmp3747[139], tmp3747[138], tmp3747[137], tmp3747[136], tmp3747[135], tmp3747[134], tmp3747[133], tmp3747[132], tmp3747[131], tmp3747[130], tmp3747[129], tmp3747[128], tmp3747[127], tmp3747[126], tmp3747[125], tmp3747[124], tmp3747[123], tmp3747[122], tmp3747[121], tmp3747[120], tmp3747[119], tmp3747[118], tmp3747[117], tmp3747[116], tmp3747[115], tmp3747[114], tmp3747[113], tmp3747[112], tmp3747[111], tmp3747[110], tmp3747[109], tmp3747[108], tmp3747[107], tmp3747[106], tmp3747[105], tmp3747[104], tmp3747[103], tmp3747[102], tmp3747[101], tmp3747[100], tmp3747[99], tmp3747[98], tmp3747[97], tmp3747[96], tmp3747[95], tmp3747[94], tmp3747[93], tmp3747[92], tmp3747[91], tmp3747[90], tmp3747[89], tmp3747[88], tmp3747[87], tmp3747[86], tmp3747[85], tmp3747[84], tmp3747[83], tmp3747[82], tmp3747[81], tmp3747[80], tmp3747[79], tmp3747[78], tmp3747[77], tmp3747[76], tmp3747[75], tmp3747[74], tmp3747[73], tmp3747[72], tmp3747[71], tmp3747[70], tmp3747[69], tmp3747[68], tmp3747[67], tmp3747[66], tmp3747[65], tmp3747[64], tmp3747[63], tmp3747[62], tmp3747[61], tmp3747[60], tmp3747[59], tmp3747[58], tmp3747[57], tmp3747[56], tmp3747[55], tmp3747[54], tmp3747[53], tmp3747[52], tmp3747[51], tmp3747[50], tmp3747[49], tmp3747[48], tmp3747[47], tmp3747[46], tmp3747[45], tmp3747[44], tmp3747[43], tmp3747[42], tmp3747[41], tmp3747[40], tmp3747[39], tmp3747[38], tmp3747[37], tmp3747[36], tmp3747[35], tmp3747[34], tmp3747[33], tmp3747[32], tmp3747[31], tmp3747[30], tmp3747[29], tmp3747[28], tmp3747[27], tmp3747[26], tmp3747[25], tmp3747[24], tmp3747[23], tmp3747[22], tmp3747[21], tmp3747[20], tmp3747[19], tmp3747[18], tmp3747[17], tmp3747[16], tmp3747[15], tmp3747[14], tmp3747[13], tmp3747[12], tmp3747[11], tmp3747[10], tmp3747[9], tmp3747[8], tmp3747[7], tmp3747[6], tmp3747[5], tmp3747[4], tmp3747[3], tmp3747[2], tmp3747[1], tmp3747[0]};
    assign tmp3749 = {tmp3748[255], tmp3748[254], tmp3748[253], tmp3748[252], tmp3748[251], tmp3748[250], tmp3748[249], tmp3748[248], tmp3748[247], tmp3748[246], tmp3748[245], tmp3748[244], tmp3748[243], tmp3748[242], tmp3748[241], tmp3748[240], tmp3748[239], tmp3748[238], tmp3748[237], tmp3748[236], tmp3748[235], tmp3748[234], tmp3748[233], tmp3748[232], tmp3748[231], tmp3748[230], tmp3748[229], tmp3748[228], tmp3748[227], tmp3748[226], tmp3748[225], tmp3748[224], tmp3748[223], tmp3748[222], tmp3748[221], tmp3748[220], tmp3748[219], tmp3748[218], tmp3748[217], tmp3748[216], tmp3748[215], tmp3748[214], tmp3748[213], tmp3748[212], tmp3748[211], tmp3748[210], tmp3748[209], tmp3748[208], tmp3748[207], tmp3748[206], tmp3748[205], tmp3748[204], tmp3748[203], tmp3748[202], tmp3748[201], tmp3748[200], tmp3748[199], tmp3748[198], tmp3748[197], tmp3748[196], tmp3748[195], tmp3748[194], tmp3748[193], tmp3748[192], tmp3748[191], tmp3748[190], tmp3748[189], tmp3748[188], tmp3748[187], tmp3748[186], tmp3748[185], tmp3748[184], tmp3748[183], tmp3748[182], tmp3748[181], tmp3748[180], tmp3748[179], tmp3748[178], tmp3748[177], tmp3748[176], tmp3748[175], tmp3748[174], tmp3748[173], tmp3748[172], tmp3748[171], tmp3748[170], tmp3748[169], tmp3748[168], tmp3748[167], tmp3748[166], tmp3748[165], tmp3748[164], tmp3748[163], tmp3748[162], tmp3748[161], tmp3748[160], tmp3748[159], tmp3748[158], tmp3748[157], tmp3748[156], tmp3748[155], tmp3748[154], tmp3748[153], tmp3748[152], tmp3748[151], tmp3748[150], tmp3748[149], tmp3748[148], tmp3748[147], tmp3748[146], tmp3748[145], tmp3748[144], tmp3748[143], tmp3748[142], tmp3748[141], tmp3748[140], tmp3748[139], tmp3748[138], tmp3748[137], tmp3748[136], tmp3748[135], tmp3748[134], tmp3748[133], tmp3748[132], tmp3748[131], tmp3748[130], tmp3748[129], tmp3748[128], tmp3748[127], tmp3748[126], tmp3748[125], tmp3748[124], tmp3748[123], tmp3748[122], tmp3748[121], tmp3748[120], tmp3748[119], tmp3748[118], tmp3748[117], tmp3748[116], tmp3748[115], tmp3748[114], tmp3748[113], tmp3748[112], tmp3748[111], tmp3748[110], tmp3748[109], tmp3748[108], tmp3748[107], tmp3748[106], tmp3748[105], tmp3748[104], tmp3748[103], tmp3748[102], tmp3748[101], tmp3748[100], tmp3748[99], tmp3748[98], tmp3748[97], tmp3748[96], tmp3748[95], tmp3748[94], tmp3748[93], tmp3748[92], tmp3748[91], tmp3748[90], tmp3748[89], tmp3748[88], tmp3748[87], tmp3748[86], tmp3748[85], tmp3748[84], tmp3748[83], tmp3748[82], tmp3748[81], tmp3748[80], tmp3748[79], tmp3748[78], tmp3748[77], tmp3748[76], tmp3748[75], tmp3748[74], tmp3748[73], tmp3748[72], tmp3748[71], tmp3748[70], tmp3748[69], tmp3748[68], tmp3748[67], tmp3748[66], tmp3748[65], tmp3748[64], tmp3748[63], tmp3748[62], tmp3748[61], tmp3748[60], tmp3748[59], tmp3748[58], tmp3748[57], tmp3748[56], tmp3748[55], tmp3748[54], tmp3748[53], tmp3748[52], tmp3748[51], tmp3748[50], tmp3748[49], tmp3748[48], tmp3748[47], tmp3748[46], tmp3748[45], tmp3748[44], tmp3748[43], tmp3748[42], tmp3748[41], tmp3748[40], tmp3748[39], tmp3748[38], tmp3748[37], tmp3748[36], tmp3748[35], tmp3748[34], tmp3748[33], tmp3748[32], tmp3748[31], tmp3748[30], tmp3748[29], tmp3748[28], tmp3748[27], tmp3748[26], tmp3748[25], tmp3748[24], tmp3748[23], tmp3748[22], tmp3748[21], tmp3748[20], tmp3748[19], tmp3748[18], tmp3748[17], tmp3748[16], tmp3748[15], tmp3748[14], tmp3748[13], tmp3748[12], tmp3748[11], tmp3748[10], tmp3748[9], tmp3748[8], tmp3748[7], tmp3748[6], tmp3748[5], tmp3748[4], tmp3748[3], tmp3748[2], tmp3748[1], tmp3748[0]};
    assign tmp3750 = {const_380_0};
    assign tmp3751 = {tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750, tmp3750};
    assign tmp3752 = {tmp3751, const_380_0};
    assign tmp3753 = {tmp27[255]};
    assign tmp3754 = tmp3752 - tmp27;
    assign tmp3755 = {tmp3754[256]};
    assign tmp3756 = {tmp3752[255]};
    assign tmp3757 = ~tmp3756;
    assign tmp3758 = tmp3755 ^ tmp3757;
    assign tmp3759 = {tmp27[255]};
    assign tmp3760 = ~tmp3759;
    assign tmp3761 = tmp3758 ^ tmp3760;
    assign tmp3762 = {const_381_0};
    assign tmp3763 = {tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762, tmp3762};
    assign tmp3764 = {tmp3763, const_381_0};
    assign tmp3765 = {tmp3740[256]};
    assign tmp3766 = tmp3764 - tmp3740;
    assign tmp3767 = {tmp3766[257]};
    assign tmp3768 = {tmp3764[256]};
    assign tmp3769 = ~tmp3768;
    assign tmp3770 = tmp3767 ^ tmp3769;
    assign tmp3771 = {tmp3740[256]};
    assign tmp3772 = ~tmp3771;
    assign tmp3773 = tmp3770 ^ tmp3772;
    assign tmp3774 = tmp3761 & tmp3773;
    assign tmp3775 = {tmp3749[255]};
    assign tmp3776 = {const_382_0};
    assign tmp3777 = {tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776, tmp3776};
    assign tmp3778 = {tmp3777, const_382_0};
    assign tmp3779 = tmp3749 - tmp3778;
    assign tmp3780 = {tmp3779[256]};
    assign tmp3781 = {tmp3749[255]};
    assign tmp3782 = ~tmp3781;
    assign tmp3783 = tmp3780 ^ tmp3782;
    assign tmp3784 = {tmp3778[255]};
    assign tmp3785 = ~tmp3784;
    assign tmp3786 = tmp3783 ^ tmp3785;
    assign tmp3787 = tmp3749 == tmp3778;
    assign tmp3788 = tmp3786 | tmp3787;
    assign tmp3789 = tmp3774 & tmp3788;
    assign tmp3790 = {tmp27[255]};
    assign tmp3791 = {const_383_0};
    assign tmp3792 = {tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791, tmp3791};
    assign tmp3793 = {tmp3792, const_383_0};
    assign tmp3794 = tmp27 - tmp3793;
    assign tmp3795 = {tmp3794[256]};
    assign tmp3796 = {tmp27[255]};
    assign tmp3797 = ~tmp3796;
    assign tmp3798 = tmp3795 ^ tmp3797;
    assign tmp3799 = {tmp3793[255]};
    assign tmp3800 = ~tmp3799;
    assign tmp3801 = tmp3798 ^ tmp3800;
    assign tmp3802 = {tmp3740[256]};
    assign tmp3803 = {const_384_0};
    assign tmp3804 = {tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803, tmp3803};
    assign tmp3805 = {tmp3804, const_384_0};
    assign tmp3806 = tmp3740 - tmp3805;
    assign tmp3807 = {tmp3806[257]};
    assign tmp3808 = {tmp3740[256]};
    assign tmp3809 = ~tmp3808;
    assign tmp3810 = tmp3807 ^ tmp3809;
    assign tmp3811 = {tmp3805[256]};
    assign tmp3812 = ~tmp3811;
    assign tmp3813 = tmp3810 ^ tmp3812;
    assign tmp3814 = tmp3801 & tmp3813;
    assign tmp3815 = {const_385_0};
    assign tmp3816 = {tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815, tmp3815};
    assign tmp3817 = {tmp3816, const_385_0};
    assign tmp3818 = {tmp3749[255]};
    assign tmp3819 = tmp3817 - tmp3749;
    assign tmp3820 = {tmp3819[256]};
    assign tmp3821 = {tmp3817[255]};
    assign tmp3822 = ~tmp3821;
    assign tmp3823 = tmp3820 ^ tmp3822;
    assign tmp3824 = {tmp3749[255]};
    assign tmp3825 = ~tmp3824;
    assign tmp3826 = tmp3823 ^ tmp3825;
    assign tmp3827 = tmp3817 == tmp3749;
    assign tmp3828 = tmp3826 | tmp3827;
    assign tmp3829 = tmp3814 & tmp3828;
    assign tmp3830 = tmp3789 ? const_386_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp3749;
    assign tmp3831 = tmp3829 ? _ver_out_tmp_84 : tmp3830;
    assign tmp3832 = ~tmp35;
    assign tmp3833 = ~tmp36;
    assign tmp3834 = tmp3832 & tmp3833;
    assign tmp3835 = ~tmp57;
    assign tmp3836 = tmp3834 & tmp3835;
    assign tmp3837 = ~tmp1034;
    assign tmp3838 = tmp3836 & tmp3837;
    assign tmp3839 = tmp3838 & tmp2071;
    assign tmp3840 = ~tmp2583;
    assign tmp3841 = tmp3839 & tmp3840;
    assign tmp3842 = tmp3841 & tmp23;
    assign tmp3843 = ~tmp2627;
    assign tmp3844 = tmp3842 & tmp3843;
    assign tmp3845 = ~tmp2798;
    assign tmp3846 = tmp3844 & tmp3845;
    assign tmp3847 = tmp3846 & tmp3425;
    assign tmp3848 = ~tmp35;
    assign tmp3849 = ~tmp36;
    assign tmp3850 = tmp3848 & tmp3849;
    assign tmp3851 = ~tmp57;
    assign tmp3852 = tmp3850 & tmp3851;
    assign tmp3853 = ~tmp1034;
    assign tmp3854 = tmp3852 & tmp3853;
    assign tmp3855 = tmp3854 & tmp2071;
    assign tmp3856 = ~tmp2583;
    assign tmp3857 = tmp3855 & tmp3856;
    assign tmp3858 = tmp3857 & tmp23;
    assign tmp3859 = ~tmp2627;
    assign tmp3860 = tmp3858 & tmp3859;
    assign tmp3861 = ~tmp2798;
    assign tmp3862 = tmp3860 & tmp3861;
    assign tmp3863 = tmp3862 & tmp3425;
    assign tmp3864 = _ver_out_tmp_85 == tmp32;
    assign tmp3865 = {const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0, const_390_0};
    assign tmp3866 = {tmp3865, const_389_0};
    assign tmp3867 = tmp3866 - tmp32;
    assign tmp3868 = {const_392_0, const_392_0};
    assign tmp3869 = {tmp3868, const_391_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp3870 = tmp3864 ? tmp3869 : tmp3867;
    assign tmp3871 = {tmp28[255]};
    assign tmp3872 = {tmp3871, tmp3871};
    assign tmp3873 = {tmp3872, tmp28};
    assign tmp3874 = {tmp3870[256]};
    assign tmp3875 = {tmp3874};
    assign tmp3876 = {tmp3875, tmp3870};
    assign tmp3877 = tmp3873 + tmp3876;
    assign tmp3878 = {tmp3877[257], tmp3877[256], tmp3877[255], tmp3877[254], tmp3877[253], tmp3877[252], tmp3877[251], tmp3877[250], tmp3877[249], tmp3877[248], tmp3877[247], tmp3877[246], tmp3877[245], tmp3877[244], tmp3877[243], tmp3877[242], tmp3877[241], tmp3877[240], tmp3877[239], tmp3877[238], tmp3877[237], tmp3877[236], tmp3877[235], tmp3877[234], tmp3877[233], tmp3877[232], tmp3877[231], tmp3877[230], tmp3877[229], tmp3877[228], tmp3877[227], tmp3877[226], tmp3877[225], tmp3877[224], tmp3877[223], tmp3877[222], tmp3877[221], tmp3877[220], tmp3877[219], tmp3877[218], tmp3877[217], tmp3877[216], tmp3877[215], tmp3877[214], tmp3877[213], tmp3877[212], tmp3877[211], tmp3877[210], tmp3877[209], tmp3877[208], tmp3877[207], tmp3877[206], tmp3877[205], tmp3877[204], tmp3877[203], tmp3877[202], tmp3877[201], tmp3877[200], tmp3877[199], tmp3877[198], tmp3877[197], tmp3877[196], tmp3877[195], tmp3877[194], tmp3877[193], tmp3877[192], tmp3877[191], tmp3877[190], tmp3877[189], tmp3877[188], tmp3877[187], tmp3877[186], tmp3877[185], tmp3877[184], tmp3877[183], tmp3877[182], tmp3877[181], tmp3877[180], tmp3877[179], tmp3877[178], tmp3877[177], tmp3877[176], tmp3877[175], tmp3877[174], tmp3877[173], tmp3877[172], tmp3877[171], tmp3877[170], tmp3877[169], tmp3877[168], tmp3877[167], tmp3877[166], tmp3877[165], tmp3877[164], tmp3877[163], tmp3877[162], tmp3877[161], tmp3877[160], tmp3877[159], tmp3877[158], tmp3877[157], tmp3877[156], tmp3877[155], tmp3877[154], tmp3877[153], tmp3877[152], tmp3877[151], tmp3877[150], tmp3877[149], tmp3877[148], tmp3877[147], tmp3877[146], tmp3877[145], tmp3877[144], tmp3877[143], tmp3877[142], tmp3877[141], tmp3877[140], tmp3877[139], tmp3877[138], tmp3877[137], tmp3877[136], tmp3877[135], tmp3877[134], tmp3877[133], tmp3877[132], tmp3877[131], tmp3877[130], tmp3877[129], tmp3877[128], tmp3877[127], tmp3877[126], tmp3877[125], tmp3877[124], tmp3877[123], tmp3877[122], tmp3877[121], tmp3877[120], tmp3877[119], tmp3877[118], tmp3877[117], tmp3877[116], tmp3877[115], tmp3877[114], tmp3877[113], tmp3877[112], tmp3877[111], tmp3877[110], tmp3877[109], tmp3877[108], tmp3877[107], tmp3877[106], tmp3877[105], tmp3877[104], tmp3877[103], tmp3877[102], tmp3877[101], tmp3877[100], tmp3877[99], tmp3877[98], tmp3877[97], tmp3877[96], tmp3877[95], tmp3877[94], tmp3877[93], tmp3877[92], tmp3877[91], tmp3877[90], tmp3877[89], tmp3877[88], tmp3877[87], tmp3877[86], tmp3877[85], tmp3877[84], tmp3877[83], tmp3877[82], tmp3877[81], tmp3877[80], tmp3877[79], tmp3877[78], tmp3877[77], tmp3877[76], tmp3877[75], tmp3877[74], tmp3877[73], tmp3877[72], tmp3877[71], tmp3877[70], tmp3877[69], tmp3877[68], tmp3877[67], tmp3877[66], tmp3877[65], tmp3877[64], tmp3877[63], tmp3877[62], tmp3877[61], tmp3877[60], tmp3877[59], tmp3877[58], tmp3877[57], tmp3877[56], tmp3877[55], tmp3877[54], tmp3877[53], tmp3877[52], tmp3877[51], tmp3877[50], tmp3877[49], tmp3877[48], tmp3877[47], tmp3877[46], tmp3877[45], tmp3877[44], tmp3877[43], tmp3877[42], tmp3877[41], tmp3877[40], tmp3877[39], tmp3877[38], tmp3877[37], tmp3877[36], tmp3877[35], tmp3877[34], tmp3877[33], tmp3877[32], tmp3877[31], tmp3877[30], tmp3877[29], tmp3877[28], tmp3877[27], tmp3877[26], tmp3877[25], tmp3877[24], tmp3877[23], tmp3877[22], tmp3877[21], tmp3877[20], tmp3877[19], tmp3877[18], tmp3877[17], tmp3877[16], tmp3877[15], tmp3877[14], tmp3877[13], tmp3877[12], tmp3877[11], tmp3877[10], tmp3877[9], tmp3877[8], tmp3877[7], tmp3877[6], tmp3877[5], tmp3877[4], tmp3877[3], tmp3877[2], tmp3877[1], tmp3877[0]};
    assign tmp3879 = {tmp3878[255], tmp3878[254], tmp3878[253], tmp3878[252], tmp3878[251], tmp3878[250], tmp3878[249], tmp3878[248], tmp3878[247], tmp3878[246], tmp3878[245], tmp3878[244], tmp3878[243], tmp3878[242], tmp3878[241], tmp3878[240], tmp3878[239], tmp3878[238], tmp3878[237], tmp3878[236], tmp3878[235], tmp3878[234], tmp3878[233], tmp3878[232], tmp3878[231], tmp3878[230], tmp3878[229], tmp3878[228], tmp3878[227], tmp3878[226], tmp3878[225], tmp3878[224], tmp3878[223], tmp3878[222], tmp3878[221], tmp3878[220], tmp3878[219], tmp3878[218], tmp3878[217], tmp3878[216], tmp3878[215], tmp3878[214], tmp3878[213], tmp3878[212], tmp3878[211], tmp3878[210], tmp3878[209], tmp3878[208], tmp3878[207], tmp3878[206], tmp3878[205], tmp3878[204], tmp3878[203], tmp3878[202], tmp3878[201], tmp3878[200], tmp3878[199], tmp3878[198], tmp3878[197], tmp3878[196], tmp3878[195], tmp3878[194], tmp3878[193], tmp3878[192], tmp3878[191], tmp3878[190], tmp3878[189], tmp3878[188], tmp3878[187], tmp3878[186], tmp3878[185], tmp3878[184], tmp3878[183], tmp3878[182], tmp3878[181], tmp3878[180], tmp3878[179], tmp3878[178], tmp3878[177], tmp3878[176], tmp3878[175], tmp3878[174], tmp3878[173], tmp3878[172], tmp3878[171], tmp3878[170], tmp3878[169], tmp3878[168], tmp3878[167], tmp3878[166], tmp3878[165], tmp3878[164], tmp3878[163], tmp3878[162], tmp3878[161], tmp3878[160], tmp3878[159], tmp3878[158], tmp3878[157], tmp3878[156], tmp3878[155], tmp3878[154], tmp3878[153], tmp3878[152], tmp3878[151], tmp3878[150], tmp3878[149], tmp3878[148], tmp3878[147], tmp3878[146], tmp3878[145], tmp3878[144], tmp3878[143], tmp3878[142], tmp3878[141], tmp3878[140], tmp3878[139], tmp3878[138], tmp3878[137], tmp3878[136], tmp3878[135], tmp3878[134], tmp3878[133], tmp3878[132], tmp3878[131], tmp3878[130], tmp3878[129], tmp3878[128], tmp3878[127], tmp3878[126], tmp3878[125], tmp3878[124], tmp3878[123], tmp3878[122], tmp3878[121], tmp3878[120], tmp3878[119], tmp3878[118], tmp3878[117], tmp3878[116], tmp3878[115], tmp3878[114], tmp3878[113], tmp3878[112], tmp3878[111], tmp3878[110], tmp3878[109], tmp3878[108], tmp3878[107], tmp3878[106], tmp3878[105], tmp3878[104], tmp3878[103], tmp3878[102], tmp3878[101], tmp3878[100], tmp3878[99], tmp3878[98], tmp3878[97], tmp3878[96], tmp3878[95], tmp3878[94], tmp3878[93], tmp3878[92], tmp3878[91], tmp3878[90], tmp3878[89], tmp3878[88], tmp3878[87], tmp3878[86], tmp3878[85], tmp3878[84], tmp3878[83], tmp3878[82], tmp3878[81], tmp3878[80], tmp3878[79], tmp3878[78], tmp3878[77], tmp3878[76], tmp3878[75], tmp3878[74], tmp3878[73], tmp3878[72], tmp3878[71], tmp3878[70], tmp3878[69], tmp3878[68], tmp3878[67], tmp3878[66], tmp3878[65], tmp3878[64], tmp3878[63], tmp3878[62], tmp3878[61], tmp3878[60], tmp3878[59], tmp3878[58], tmp3878[57], tmp3878[56], tmp3878[55], tmp3878[54], tmp3878[53], tmp3878[52], tmp3878[51], tmp3878[50], tmp3878[49], tmp3878[48], tmp3878[47], tmp3878[46], tmp3878[45], tmp3878[44], tmp3878[43], tmp3878[42], tmp3878[41], tmp3878[40], tmp3878[39], tmp3878[38], tmp3878[37], tmp3878[36], tmp3878[35], tmp3878[34], tmp3878[33], tmp3878[32], tmp3878[31], tmp3878[30], tmp3878[29], tmp3878[28], tmp3878[27], tmp3878[26], tmp3878[25], tmp3878[24], tmp3878[23], tmp3878[22], tmp3878[21], tmp3878[20], tmp3878[19], tmp3878[18], tmp3878[17], tmp3878[16], tmp3878[15], tmp3878[14], tmp3878[13], tmp3878[12], tmp3878[11], tmp3878[10], tmp3878[9], tmp3878[8], tmp3878[7], tmp3878[6], tmp3878[5], tmp3878[4], tmp3878[3], tmp3878[2], tmp3878[1], tmp3878[0]};
    assign tmp3880 = {const_393_0};
    assign tmp3881 = {tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880, tmp3880};
    assign tmp3882 = {tmp3881, const_393_0};
    assign tmp3883 = {tmp28[255]};
    assign tmp3884 = tmp3882 - tmp28;
    assign tmp3885 = {tmp3884[256]};
    assign tmp3886 = {tmp3882[255]};
    assign tmp3887 = ~tmp3886;
    assign tmp3888 = tmp3885 ^ tmp3887;
    assign tmp3889 = {tmp28[255]};
    assign tmp3890 = ~tmp3889;
    assign tmp3891 = tmp3888 ^ tmp3890;
    assign tmp3892 = {const_394_0};
    assign tmp3893 = {tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892, tmp3892};
    assign tmp3894 = {tmp3893, const_394_0};
    assign tmp3895 = {tmp3870[256]};
    assign tmp3896 = tmp3894 - tmp3870;
    assign tmp3897 = {tmp3896[257]};
    assign tmp3898 = {tmp3894[256]};
    assign tmp3899 = ~tmp3898;
    assign tmp3900 = tmp3897 ^ tmp3899;
    assign tmp3901 = {tmp3870[256]};
    assign tmp3902 = ~tmp3901;
    assign tmp3903 = tmp3900 ^ tmp3902;
    assign tmp3904 = tmp3891 & tmp3903;
    assign tmp3905 = {tmp3879[255]};
    assign tmp3906 = {const_395_0};
    assign tmp3907 = {tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906, tmp3906};
    assign tmp3908 = {tmp3907, const_395_0};
    assign tmp3909 = tmp3879 - tmp3908;
    assign tmp3910 = {tmp3909[256]};
    assign tmp3911 = {tmp3879[255]};
    assign tmp3912 = ~tmp3911;
    assign tmp3913 = tmp3910 ^ tmp3912;
    assign tmp3914 = {tmp3908[255]};
    assign tmp3915 = ~tmp3914;
    assign tmp3916 = tmp3913 ^ tmp3915;
    assign tmp3917 = tmp3879 == tmp3908;
    assign tmp3918 = tmp3916 | tmp3917;
    assign tmp3919 = tmp3904 & tmp3918;
    assign tmp3920 = {tmp28[255]};
    assign tmp3921 = {const_396_0};
    assign tmp3922 = {tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921, tmp3921};
    assign tmp3923 = {tmp3922, const_396_0};
    assign tmp3924 = tmp28 - tmp3923;
    assign tmp3925 = {tmp3924[256]};
    assign tmp3926 = {tmp28[255]};
    assign tmp3927 = ~tmp3926;
    assign tmp3928 = tmp3925 ^ tmp3927;
    assign tmp3929 = {tmp3923[255]};
    assign tmp3930 = ~tmp3929;
    assign tmp3931 = tmp3928 ^ tmp3930;
    assign tmp3932 = {tmp3870[256]};
    assign tmp3933 = {const_397_0};
    assign tmp3934 = {tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933, tmp3933};
    assign tmp3935 = {tmp3934, const_397_0};
    assign tmp3936 = tmp3870 - tmp3935;
    assign tmp3937 = {tmp3936[257]};
    assign tmp3938 = {tmp3870[256]};
    assign tmp3939 = ~tmp3938;
    assign tmp3940 = tmp3937 ^ tmp3939;
    assign tmp3941 = {tmp3935[256]};
    assign tmp3942 = ~tmp3941;
    assign tmp3943 = tmp3940 ^ tmp3942;
    assign tmp3944 = tmp3931 & tmp3943;
    assign tmp3945 = {const_398_0};
    assign tmp3946 = {tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945, tmp3945};
    assign tmp3947 = {tmp3946, const_398_0};
    assign tmp3948 = {tmp3879[255]};
    assign tmp3949 = tmp3947 - tmp3879;
    assign tmp3950 = {tmp3949[256]};
    assign tmp3951 = {tmp3947[255]};
    assign tmp3952 = ~tmp3951;
    assign tmp3953 = tmp3950 ^ tmp3952;
    assign tmp3954 = {tmp3879[255]};
    assign tmp3955 = ~tmp3954;
    assign tmp3956 = tmp3953 ^ tmp3955;
    assign tmp3957 = tmp3947 == tmp3879;
    assign tmp3958 = tmp3956 | tmp3957;
    assign tmp3959 = tmp3944 & tmp3958;
    assign tmp3960 = tmp3919 ? const_399_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp3879;
    assign tmp3961 = tmp3959 ? _ver_out_tmp_87 : tmp3960;
    assign tmp3962 = ~tmp35;
    assign tmp3963 = ~tmp36;
    assign tmp3964 = tmp3962 & tmp3963;
    assign tmp3965 = ~tmp57;
    assign tmp3966 = tmp3964 & tmp3965;
    assign tmp3967 = ~tmp1034;
    assign tmp3968 = tmp3966 & tmp3967;
    assign tmp3969 = tmp3968 & tmp2071;
    assign tmp3970 = ~tmp2583;
    assign tmp3971 = tmp3969 & tmp3970;
    assign tmp3972 = tmp3971 & tmp23;
    assign tmp3973 = ~tmp2627;
    assign tmp3974 = tmp3972 & tmp3973;
    assign tmp3975 = ~tmp2798;
    assign tmp3976 = tmp3974 & tmp3975;
    assign tmp3977 = tmp3976 & tmp3425;
    assign tmp3978 = {tmp25[255]};
    assign tmp3979 = {tmp29[255]};
    assign tmp3980 = tmp25 - tmp29;
    assign tmp3981 = {tmp3980[256]};
    assign tmp3982 = {tmp25[255]};
    assign tmp3983 = ~tmp3982;
    assign tmp3984 = tmp3981 ^ tmp3983;
    assign tmp3985 = {tmp29[255]};
    assign tmp3986 = ~tmp3985;
    assign tmp3987 = tmp3984 ^ tmp3986;
    assign tmp3988 = {tmp26[255]};
    assign tmp3989 = {tmp30[255]};
    assign tmp3990 = tmp26 - tmp30;
    assign tmp3991 = {tmp3990[256]};
    assign tmp3992 = {tmp26[255]};
    assign tmp3993 = ~tmp3992;
    assign tmp3994 = tmp3991 ^ tmp3993;
    assign tmp3995 = {tmp30[255]};
    assign tmp3996 = ~tmp3995;
    assign tmp3997 = tmp3994 ^ tmp3996;
    assign tmp3998 = tmp3987 & tmp3997;
    assign tmp3999 = {tmp27[255]};
    assign tmp4000 = {tmp31[255]};
    assign tmp4001 = tmp27 - tmp31;
    assign tmp4002 = {tmp4001[256]};
    assign tmp4003 = {tmp27[255]};
    assign tmp4004 = ~tmp4003;
    assign tmp4005 = tmp4002 ^ tmp4004;
    assign tmp4006 = {tmp31[255]};
    assign tmp4007 = ~tmp4006;
    assign tmp4008 = tmp4005 ^ tmp4007;
    assign tmp4009 = tmp3998 & tmp4008;
    assign tmp4010 = {tmp28[255]};
    assign tmp4011 = {tmp32[255]};
    assign tmp4012 = tmp28 - tmp32;
    assign tmp4013 = {tmp4012[256]};
    assign tmp4014 = {tmp28[255]};
    assign tmp4015 = ~tmp4014;
    assign tmp4016 = tmp4013 ^ tmp4015;
    assign tmp4017 = {tmp32[255]};
    assign tmp4018 = ~tmp4017;
    assign tmp4019 = tmp4016 ^ tmp4018;
    assign tmp4020 = tmp4009 & tmp4019;
    assign tmp4021 = ~tmp35;
    assign tmp4022 = ~tmp36;
    assign tmp4023 = tmp4021 & tmp4022;
    assign tmp4024 = ~tmp57;
    assign tmp4025 = tmp4023 & tmp4024;
    assign tmp4026 = ~tmp1034;
    assign tmp4027 = tmp4025 & tmp4026;
    assign tmp4028 = tmp4027 & tmp2071;
    assign tmp4029 = ~tmp2583;
    assign tmp4030 = tmp4028 & tmp4029;
    assign tmp4031 = tmp4030 & tmp23;
    assign tmp4032 = ~tmp2627;
    assign tmp4033 = tmp4031 & tmp4032;
    assign tmp4034 = ~tmp2798;
    assign tmp4035 = tmp4033 & tmp4034;
    assign tmp4036 = ~tmp3425;
    assign tmp4037 = tmp4035 & tmp4036;
    assign tmp4038 = tmp4037 & tmp4020;
    assign tmp4039 = ~tmp35;
    assign tmp4040 = ~tmp36;
    assign tmp4041 = tmp4039 & tmp4040;
    assign tmp4042 = ~tmp57;
    assign tmp4043 = tmp4041 & tmp4042;
    assign tmp4044 = ~tmp1034;
    assign tmp4045 = tmp4043 & tmp4044;
    assign tmp4046 = tmp4045 & tmp2071;
    assign tmp4047 = ~tmp2583;
    assign tmp4048 = tmp4046 & tmp4047;
    assign tmp4049 = tmp4048 & tmp23;
    assign tmp4050 = ~tmp2627;
    assign tmp4051 = tmp4049 & tmp4050;
    assign tmp4052 = ~tmp2798;
    assign tmp4053 = tmp4051 & tmp4052;
    assign tmp4054 = ~tmp3425;
    assign tmp4055 = tmp4053 & tmp4054;
    assign tmp4056 = tmp4055 & tmp4020;
    assign tmp4057 = ~tmp35;
    assign tmp4058 = ~tmp36;
    assign tmp4059 = tmp4057 & tmp4058;
    assign tmp4060 = ~tmp57;
    assign tmp4061 = tmp4059 & tmp4060;
    assign tmp4062 = ~tmp1034;
    assign tmp4063 = tmp4061 & tmp4062;
    assign tmp4064 = tmp4063 & tmp2071;
    assign tmp4065 = ~tmp2583;
    assign tmp4066 = tmp4064 & tmp4065;
    assign tmp4067 = tmp4066 & tmp23;
    assign tmp4068 = ~tmp2627;
    assign tmp4069 = tmp4067 & tmp4068;
    assign tmp4070 = ~tmp2798;
    assign tmp4071 = tmp4069 & tmp4070;
    assign tmp4072 = ~tmp3425;
    assign tmp4073 = tmp4071 & tmp4072;
    assign tmp4074 = tmp4073 & tmp4020;
    assign tmp4075 = ~tmp35;
    assign tmp4076 = ~tmp36;
    assign tmp4077 = tmp4075 & tmp4076;
    assign tmp4078 = ~tmp57;
    assign tmp4079 = tmp4077 & tmp4078;
    assign tmp4080 = ~tmp1034;
    assign tmp4081 = tmp4079 & tmp4080;
    assign tmp4082 = tmp4081 & tmp2071;
    assign tmp4083 = ~tmp2583;
    assign tmp4084 = tmp4082 & tmp4083;
    assign tmp4085 = tmp4084 & tmp23;
    assign tmp4086 = ~tmp2627;
    assign tmp4087 = tmp4085 & tmp4086;
    assign tmp4088 = ~tmp2798;
    assign tmp4089 = tmp4087 & tmp4088;
    assign tmp4090 = ~tmp3425;
    assign tmp4091 = tmp4089 & tmp4090;
    assign tmp4092 = tmp4091 & tmp4020;
    assign tmp4093 = ~tmp35;
    assign tmp4094 = ~tmp36;
    assign tmp4095 = tmp4093 & tmp4094;
    assign tmp4096 = ~tmp57;
    assign tmp4097 = tmp4095 & tmp4096;
    assign tmp4098 = ~tmp1034;
    assign tmp4099 = tmp4097 & tmp4098;
    assign tmp4100 = tmp4099 & tmp2071;
    assign tmp4101 = ~tmp2583;
    assign tmp4102 = tmp4100 & tmp4101;
    assign tmp4103 = tmp4102 & tmp23;
    assign tmp4104 = ~tmp2627;
    assign tmp4105 = tmp4103 & tmp4104;
    assign tmp4106 = ~tmp2798;
    assign tmp4107 = tmp4105 & tmp4106;
    assign tmp4108 = ~tmp3425;
    assign tmp4109 = tmp4107 & tmp4108;
    assign tmp4110 = tmp4109 & tmp4020;
    assign tmp4111 = ~tmp35;
    assign tmp4112 = ~tmp36;
    assign tmp4113 = tmp4111 & tmp4112;
    assign tmp4114 = ~tmp57;
    assign tmp4115 = tmp4113 & tmp4114;
    assign tmp4116 = ~tmp1034;
    assign tmp4117 = tmp4115 & tmp4116;
    assign tmp4118 = tmp4117 & tmp2071;
    assign tmp4119 = ~tmp2583;
    assign tmp4120 = tmp4118 & tmp4119;
    assign tmp4121 = tmp4120 & tmp23;
    assign tmp4122 = ~tmp2627;
    assign tmp4123 = tmp4121 & tmp4122;
    assign tmp4124 = ~tmp2798;
    assign tmp4125 = tmp4123 & tmp4124;
    assign tmp4126 = ~tmp3425;
    assign tmp4127 = tmp4125 & tmp4126;
    assign tmp4128 = tmp4127 & tmp4020;
    assign tmp4129 = ~tmp35;
    assign tmp4130 = ~tmp36;
    assign tmp4131 = tmp4129 & tmp4130;
    assign tmp4132 = ~tmp57;
    assign tmp4133 = tmp4131 & tmp4132;
    assign tmp4134 = ~tmp1034;
    assign tmp4135 = tmp4133 & tmp4134;
    assign tmp4136 = tmp4135 & tmp2071;
    assign tmp4137 = ~tmp2583;
    assign tmp4138 = tmp4136 & tmp4137;
    assign tmp4139 = tmp4138 & tmp23;
    assign tmp4140 = ~tmp2627;
    assign tmp4141 = tmp4139 & tmp4140;
    assign tmp4142 = ~tmp2798;
    assign tmp4143 = tmp4141 & tmp4142;
    assign tmp4144 = ~tmp3425;
    assign tmp4145 = tmp4143 & tmp4144;
    assign tmp4146 = tmp4145 & tmp4020;
    assign tmp4147 = ~tmp35;
    assign tmp4148 = ~tmp36;
    assign tmp4149 = tmp4147 & tmp4148;
    assign tmp4150 = ~tmp57;
    assign tmp4151 = tmp4149 & tmp4150;
    assign tmp4152 = ~tmp1034;
    assign tmp4153 = tmp4151 & tmp4152;
    assign tmp4154 = tmp4153 & tmp2071;
    assign tmp4155 = ~tmp2583;
    assign tmp4156 = tmp4154 & tmp4155;
    assign tmp4157 = tmp4156 & tmp23;
    assign tmp4158 = ~tmp2627;
    assign tmp4159 = tmp4157 & tmp4158;
    assign tmp4160 = ~tmp2798;
    assign tmp4161 = tmp4159 & tmp4160;
    assign tmp4162 = ~tmp3425;
    assign tmp4163 = tmp4161 & tmp4162;
    assign tmp4164 = tmp4163 & tmp4020;
    assign tmp4165 = ~tmp35;
    assign tmp4166 = ~tmp36;
    assign tmp4167 = tmp4165 & tmp4166;
    assign tmp4168 = ~tmp57;
    assign tmp4169 = tmp4167 & tmp4168;
    assign tmp4170 = ~tmp1034;
    assign tmp4171 = tmp4169 & tmp4170;
    assign tmp4172 = tmp4171 & tmp2071;
    assign tmp4173 = ~tmp2583;
    assign tmp4174 = tmp4172 & tmp4173;
    assign tmp4175 = tmp4174 & tmp23;
    assign tmp4176 = ~tmp2627;
    assign tmp4177 = tmp4175 & tmp4176;
    assign tmp4178 = ~tmp2798;
    assign tmp4179 = tmp4177 & tmp4178;
    assign tmp4180 = ~tmp3425;
    assign tmp4181 = tmp4179 & tmp4180;
    assign tmp4182 = tmp4181 & tmp4020;
    assign tmp4183 = ~tmp35;
    assign tmp4184 = ~tmp36;
    assign tmp4185 = tmp4183 & tmp4184;
    assign tmp4186 = ~tmp57;
    assign tmp4187 = tmp4185 & tmp4186;
    assign tmp4188 = ~tmp1034;
    assign tmp4189 = tmp4187 & tmp4188;
    assign tmp4190 = tmp4189 & tmp2071;
    assign tmp4191 = ~tmp2583;
    assign tmp4192 = tmp4190 & tmp4191;
    assign tmp4193 = tmp4192 & tmp23;
    assign tmp4194 = ~tmp2627;
    assign tmp4195 = tmp4193 & tmp4194;
    assign tmp4196 = ~tmp2798;
    assign tmp4197 = tmp4195 & tmp4196;
    assign tmp4198 = ~tmp3425;
    assign tmp4199 = tmp4197 & tmp4198;
    assign tmp4200 = tmp4199 & tmp4020;
    assign tmp4201 = {tmp29[255]};
    assign tmp4202 = {tmp25[255]};
    assign tmp4203 = tmp29 - tmp25;
    assign tmp4204 = {tmp4203[256]};
    assign tmp4205 = {tmp29[255]};
    assign tmp4206 = ~tmp4205;
    assign tmp4207 = tmp4204 ^ tmp4206;
    assign tmp4208 = {tmp25[255]};
    assign tmp4209 = ~tmp4208;
    assign tmp4210 = tmp4207 ^ tmp4209;
    assign tmp4211 = {tmp29[253], tmp29[252], tmp29[251], tmp29[250], tmp29[249], tmp29[248], tmp29[247], tmp29[246], tmp29[245], tmp29[244], tmp29[243], tmp29[242], tmp29[241], tmp29[240], tmp29[239], tmp29[238], tmp29[237], tmp29[236], tmp29[235], tmp29[234], tmp29[233], tmp29[232], tmp29[231], tmp29[230], tmp29[229], tmp29[228], tmp29[227], tmp29[226], tmp29[225], tmp29[224], tmp29[223], tmp29[222], tmp29[221], tmp29[220], tmp29[219], tmp29[218], tmp29[217], tmp29[216], tmp29[215], tmp29[214], tmp29[213], tmp29[212], tmp29[211], tmp29[210], tmp29[209], tmp29[208], tmp29[207], tmp29[206], tmp29[205], tmp29[204], tmp29[203], tmp29[202], tmp29[201], tmp29[200], tmp29[199], tmp29[198], tmp29[197], tmp29[196], tmp29[195], tmp29[194], tmp29[193], tmp29[192], tmp29[191], tmp29[190], tmp29[189], tmp29[188], tmp29[187], tmp29[186], tmp29[185], tmp29[184], tmp29[183], tmp29[182], tmp29[181], tmp29[180], tmp29[179], tmp29[178], tmp29[177], tmp29[176], tmp29[175], tmp29[174], tmp29[173], tmp29[172], tmp29[171], tmp29[170], tmp29[169], tmp29[168], tmp29[167], tmp29[166], tmp29[165], tmp29[164], tmp29[163], tmp29[162], tmp29[161], tmp29[160], tmp29[159], tmp29[158], tmp29[157], tmp29[156], tmp29[155], tmp29[154], tmp29[153], tmp29[152], tmp29[151], tmp29[150], tmp29[149], tmp29[148], tmp29[147], tmp29[146], tmp29[145], tmp29[144], tmp29[143], tmp29[142], tmp29[141], tmp29[140], tmp29[139], tmp29[138], tmp29[137], tmp29[136], tmp29[135], tmp29[134], tmp29[133], tmp29[132], tmp29[131], tmp29[130], tmp29[129], tmp29[128], tmp29[127], tmp29[126], tmp29[125], tmp29[124], tmp29[123], tmp29[122], tmp29[121], tmp29[120], tmp29[119], tmp29[118], tmp29[117], tmp29[116], tmp29[115], tmp29[114], tmp29[113], tmp29[112], tmp29[111], tmp29[110], tmp29[109], tmp29[108], tmp29[107], tmp29[106], tmp29[105], tmp29[104], tmp29[103], tmp29[102], tmp29[101], tmp29[100], tmp29[99], tmp29[98], tmp29[97], tmp29[96], tmp29[95], tmp29[94], tmp29[93], tmp29[92], tmp29[91], tmp29[90], tmp29[89], tmp29[88], tmp29[87], tmp29[86], tmp29[85], tmp29[84], tmp29[83], tmp29[82], tmp29[81], tmp29[80], tmp29[79], tmp29[78], tmp29[77], tmp29[76], tmp29[75], tmp29[74], tmp29[73], tmp29[72], tmp29[71], tmp29[70], tmp29[69], tmp29[68], tmp29[67], tmp29[66], tmp29[65], tmp29[64], tmp29[63], tmp29[62], tmp29[61], tmp29[60], tmp29[59], tmp29[58], tmp29[57], tmp29[56], tmp29[55], tmp29[54], tmp29[53], tmp29[52], tmp29[51], tmp29[50], tmp29[49], tmp29[48], tmp29[47], tmp29[46], tmp29[45], tmp29[44], tmp29[43], tmp29[42], tmp29[41], tmp29[40], tmp29[39], tmp29[38], tmp29[37], tmp29[36], tmp29[35], tmp29[34], tmp29[33], tmp29[32], tmp29[31], tmp29[30], tmp29[29], tmp29[28], tmp29[27], tmp29[26], tmp29[25], tmp29[24], tmp29[23], tmp29[22], tmp29[21], tmp29[20], tmp29[19], tmp29[18], tmp29[17], tmp29[16], tmp29[15], tmp29[14], tmp29[13], tmp29[12], tmp29[11], tmp29[10], tmp29[9], tmp29[8], tmp29[7], tmp29[6], tmp29[5], tmp29[4], tmp29[3], tmp29[2], tmp29[1], tmp29[0]};
    assign tmp4212 = {tmp4211, const_403_0};
    assign tmp4213 = {const_404_0};
    assign tmp4214 = {tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213, tmp4213};
    assign tmp4215 = {tmp4214, const_404_0};
    assign tmp4216 = {tmp29[255]};
    assign tmp4217 = tmp4215 - tmp29;
    assign tmp4218 = {tmp4217[256]};
    assign tmp4219 = {tmp4215[255]};
    assign tmp4220 = ~tmp4219;
    assign tmp4221 = tmp4218 ^ tmp4220;
    assign tmp4222 = {tmp29[255]};
    assign tmp4223 = ~tmp4222;
    assign tmp4224 = tmp4221 ^ tmp4223;
    assign tmp4225 = {tmp4212[255]};
    assign tmp4226 = {const_405_0};
    assign tmp4227 = {tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226, tmp4226};
    assign tmp4228 = {tmp4227, const_405_0};
    assign tmp4229 = tmp4212 - tmp4228;
    assign tmp4230 = {tmp4229[256]};
    assign tmp4231 = {tmp4212[255]};
    assign tmp4232 = ~tmp4231;
    assign tmp4233 = tmp4230 ^ tmp4232;
    assign tmp4234 = {tmp4228[255]};
    assign tmp4235 = ~tmp4234;
    assign tmp4236 = tmp4233 ^ tmp4235;
    assign tmp4237 = tmp4224 & tmp4236;
    assign tmp4238 = {tmp29[255]};
    assign tmp4239 = {const_406_0};
    assign tmp4240 = {tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239, tmp4239};
    assign tmp4241 = {tmp4240, const_406_0};
    assign tmp4242 = tmp29 - tmp4241;
    assign tmp4243 = {tmp4242[256]};
    assign tmp4244 = {tmp29[255]};
    assign tmp4245 = ~tmp4244;
    assign tmp4246 = tmp4243 ^ tmp4245;
    assign tmp4247 = {tmp4241[255]};
    assign tmp4248 = ~tmp4247;
    assign tmp4249 = tmp4246 ^ tmp4248;
    assign tmp4250 = {const_407_0};
    assign tmp4251 = {tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250, tmp4250};
    assign tmp4252 = {tmp4251, const_407_0};
    assign tmp4253 = {tmp4212[255]};
    assign tmp4254 = tmp4252 - tmp4212;
    assign tmp4255 = {tmp4254[256]};
    assign tmp4256 = {tmp4252[255]};
    assign tmp4257 = ~tmp4256;
    assign tmp4258 = tmp4255 ^ tmp4257;
    assign tmp4259 = {tmp4212[255]};
    assign tmp4260 = ~tmp4259;
    assign tmp4261 = tmp4258 ^ tmp4260;
    assign tmp4262 = tmp4252 == tmp4212;
    assign tmp4263 = tmp4261 | tmp4262;
    assign tmp4264 = tmp4249 & tmp4263;
    assign tmp4265 = tmp4237 ? const_408_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp4212;
    assign tmp4266 = tmp4264 ? _ver_out_tmp_90 : tmp4265;
    assign tmp4267 = {tmp25[255]};
    assign tmp4268 = {tmp4266[255]};
    assign tmp4269 = tmp25 - tmp4266;
    assign tmp4270 = {tmp4269[256]};
    assign tmp4271 = {tmp25[255]};
    assign tmp4272 = ~tmp4271;
    assign tmp4273 = tmp4270 ^ tmp4272;
    assign tmp4274 = {tmp4266[255]};
    assign tmp4275 = ~tmp4274;
    assign tmp4276 = tmp4273 ^ tmp4275;
    assign tmp4277 = tmp4210 & tmp4276;
    assign tmp4278 = {tmp30[255]};
    assign tmp4279 = {tmp26[255]};
    assign tmp4280 = tmp30 - tmp26;
    assign tmp4281 = {tmp4280[256]};
    assign tmp4282 = {tmp30[255]};
    assign tmp4283 = ~tmp4282;
    assign tmp4284 = tmp4281 ^ tmp4283;
    assign tmp4285 = {tmp26[255]};
    assign tmp4286 = ~tmp4285;
    assign tmp4287 = tmp4284 ^ tmp4286;
    assign tmp4288 = tmp4277 & tmp4287;
    assign tmp4289 = {tmp30[253], tmp30[252], tmp30[251], tmp30[250], tmp30[249], tmp30[248], tmp30[247], tmp30[246], tmp30[245], tmp30[244], tmp30[243], tmp30[242], tmp30[241], tmp30[240], tmp30[239], tmp30[238], tmp30[237], tmp30[236], tmp30[235], tmp30[234], tmp30[233], tmp30[232], tmp30[231], tmp30[230], tmp30[229], tmp30[228], tmp30[227], tmp30[226], tmp30[225], tmp30[224], tmp30[223], tmp30[222], tmp30[221], tmp30[220], tmp30[219], tmp30[218], tmp30[217], tmp30[216], tmp30[215], tmp30[214], tmp30[213], tmp30[212], tmp30[211], tmp30[210], tmp30[209], tmp30[208], tmp30[207], tmp30[206], tmp30[205], tmp30[204], tmp30[203], tmp30[202], tmp30[201], tmp30[200], tmp30[199], tmp30[198], tmp30[197], tmp30[196], tmp30[195], tmp30[194], tmp30[193], tmp30[192], tmp30[191], tmp30[190], tmp30[189], tmp30[188], tmp30[187], tmp30[186], tmp30[185], tmp30[184], tmp30[183], tmp30[182], tmp30[181], tmp30[180], tmp30[179], tmp30[178], tmp30[177], tmp30[176], tmp30[175], tmp30[174], tmp30[173], tmp30[172], tmp30[171], tmp30[170], tmp30[169], tmp30[168], tmp30[167], tmp30[166], tmp30[165], tmp30[164], tmp30[163], tmp30[162], tmp30[161], tmp30[160], tmp30[159], tmp30[158], tmp30[157], tmp30[156], tmp30[155], tmp30[154], tmp30[153], tmp30[152], tmp30[151], tmp30[150], tmp30[149], tmp30[148], tmp30[147], tmp30[146], tmp30[145], tmp30[144], tmp30[143], tmp30[142], tmp30[141], tmp30[140], tmp30[139], tmp30[138], tmp30[137], tmp30[136], tmp30[135], tmp30[134], tmp30[133], tmp30[132], tmp30[131], tmp30[130], tmp30[129], tmp30[128], tmp30[127], tmp30[126], tmp30[125], tmp30[124], tmp30[123], tmp30[122], tmp30[121], tmp30[120], tmp30[119], tmp30[118], tmp30[117], tmp30[116], tmp30[115], tmp30[114], tmp30[113], tmp30[112], tmp30[111], tmp30[110], tmp30[109], tmp30[108], tmp30[107], tmp30[106], tmp30[105], tmp30[104], tmp30[103], tmp30[102], tmp30[101], tmp30[100], tmp30[99], tmp30[98], tmp30[97], tmp30[96], tmp30[95], tmp30[94], tmp30[93], tmp30[92], tmp30[91], tmp30[90], tmp30[89], tmp30[88], tmp30[87], tmp30[86], tmp30[85], tmp30[84], tmp30[83], tmp30[82], tmp30[81], tmp30[80], tmp30[79], tmp30[78], tmp30[77], tmp30[76], tmp30[75], tmp30[74], tmp30[73], tmp30[72], tmp30[71], tmp30[70], tmp30[69], tmp30[68], tmp30[67], tmp30[66], tmp30[65], tmp30[64], tmp30[63], tmp30[62], tmp30[61], tmp30[60], tmp30[59], tmp30[58], tmp30[57], tmp30[56], tmp30[55], tmp30[54], tmp30[53], tmp30[52], tmp30[51], tmp30[50], tmp30[49], tmp30[48], tmp30[47], tmp30[46], tmp30[45], tmp30[44], tmp30[43], tmp30[42], tmp30[41], tmp30[40], tmp30[39], tmp30[38], tmp30[37], tmp30[36], tmp30[35], tmp30[34], tmp30[33], tmp30[32], tmp30[31], tmp30[30], tmp30[29], tmp30[28], tmp30[27], tmp30[26], tmp30[25], tmp30[24], tmp30[23], tmp30[22], tmp30[21], tmp30[20], tmp30[19], tmp30[18], tmp30[17], tmp30[16], tmp30[15], tmp30[14], tmp30[13], tmp30[12], tmp30[11], tmp30[10], tmp30[9], tmp30[8], tmp30[7], tmp30[6], tmp30[5], tmp30[4], tmp30[3], tmp30[2], tmp30[1], tmp30[0]};
    assign tmp4290 = {tmp4289, const_410_0};
    assign tmp4291 = {const_411_0};
    assign tmp4292 = {tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291, tmp4291};
    assign tmp4293 = {tmp4292, const_411_0};
    assign tmp4294 = {tmp30[255]};
    assign tmp4295 = tmp4293 - tmp30;
    assign tmp4296 = {tmp4295[256]};
    assign tmp4297 = {tmp4293[255]};
    assign tmp4298 = ~tmp4297;
    assign tmp4299 = tmp4296 ^ tmp4298;
    assign tmp4300 = {tmp30[255]};
    assign tmp4301 = ~tmp4300;
    assign tmp4302 = tmp4299 ^ tmp4301;
    assign tmp4303 = {tmp4290[255]};
    assign tmp4304 = {const_412_0};
    assign tmp4305 = {tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304, tmp4304};
    assign tmp4306 = {tmp4305, const_412_0};
    assign tmp4307 = tmp4290 - tmp4306;
    assign tmp4308 = {tmp4307[256]};
    assign tmp4309 = {tmp4290[255]};
    assign tmp4310 = ~tmp4309;
    assign tmp4311 = tmp4308 ^ tmp4310;
    assign tmp4312 = {tmp4306[255]};
    assign tmp4313 = ~tmp4312;
    assign tmp4314 = tmp4311 ^ tmp4313;
    assign tmp4315 = tmp4302 & tmp4314;
    assign tmp4316 = {tmp30[255]};
    assign tmp4317 = {const_413_0};
    assign tmp4318 = {tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317, tmp4317};
    assign tmp4319 = {tmp4318, const_413_0};
    assign tmp4320 = tmp30 - tmp4319;
    assign tmp4321 = {tmp4320[256]};
    assign tmp4322 = {tmp30[255]};
    assign tmp4323 = ~tmp4322;
    assign tmp4324 = tmp4321 ^ tmp4323;
    assign tmp4325 = {tmp4319[255]};
    assign tmp4326 = ~tmp4325;
    assign tmp4327 = tmp4324 ^ tmp4326;
    assign tmp4328 = {const_414_0};
    assign tmp4329 = {tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328, tmp4328};
    assign tmp4330 = {tmp4329, const_414_0};
    assign tmp4331 = {tmp4290[255]};
    assign tmp4332 = tmp4330 - tmp4290;
    assign tmp4333 = {tmp4332[256]};
    assign tmp4334 = {tmp4330[255]};
    assign tmp4335 = ~tmp4334;
    assign tmp4336 = tmp4333 ^ tmp4335;
    assign tmp4337 = {tmp4290[255]};
    assign tmp4338 = ~tmp4337;
    assign tmp4339 = tmp4336 ^ tmp4338;
    assign tmp4340 = tmp4330 == tmp4290;
    assign tmp4341 = tmp4339 | tmp4340;
    assign tmp4342 = tmp4327 & tmp4341;
    assign tmp4343 = tmp4315 ? const_415_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp4290;
    assign tmp4344 = tmp4342 ? _ver_out_tmp_0 : tmp4343;
    assign tmp4345 = {tmp26[255]};
    assign tmp4346 = {tmp4344[255]};
    assign tmp4347 = tmp26 - tmp4344;
    assign tmp4348 = {tmp4347[256]};
    assign tmp4349 = {tmp26[255]};
    assign tmp4350 = ~tmp4349;
    assign tmp4351 = tmp4348 ^ tmp4350;
    assign tmp4352 = {tmp4344[255]};
    assign tmp4353 = ~tmp4352;
    assign tmp4354 = tmp4351 ^ tmp4353;
    assign tmp4355 = tmp4288 & tmp4354;
    assign tmp4356 = {tmp31[255]};
    assign tmp4357 = {tmp27[255]};
    assign tmp4358 = tmp31 - tmp27;
    assign tmp4359 = {tmp4358[256]};
    assign tmp4360 = {tmp31[255]};
    assign tmp4361 = ~tmp4360;
    assign tmp4362 = tmp4359 ^ tmp4361;
    assign tmp4363 = {tmp27[255]};
    assign tmp4364 = ~tmp4363;
    assign tmp4365 = tmp4362 ^ tmp4364;
    assign tmp4366 = tmp4355 & tmp4365;
    assign tmp4367 = {tmp31[253], tmp31[252], tmp31[251], tmp31[250], tmp31[249], tmp31[248], tmp31[247], tmp31[246], tmp31[245], tmp31[244], tmp31[243], tmp31[242], tmp31[241], tmp31[240], tmp31[239], tmp31[238], tmp31[237], tmp31[236], tmp31[235], tmp31[234], tmp31[233], tmp31[232], tmp31[231], tmp31[230], tmp31[229], tmp31[228], tmp31[227], tmp31[226], tmp31[225], tmp31[224], tmp31[223], tmp31[222], tmp31[221], tmp31[220], tmp31[219], tmp31[218], tmp31[217], tmp31[216], tmp31[215], tmp31[214], tmp31[213], tmp31[212], tmp31[211], tmp31[210], tmp31[209], tmp31[208], tmp31[207], tmp31[206], tmp31[205], tmp31[204], tmp31[203], tmp31[202], tmp31[201], tmp31[200], tmp31[199], tmp31[198], tmp31[197], tmp31[196], tmp31[195], tmp31[194], tmp31[193], tmp31[192], tmp31[191], tmp31[190], tmp31[189], tmp31[188], tmp31[187], tmp31[186], tmp31[185], tmp31[184], tmp31[183], tmp31[182], tmp31[181], tmp31[180], tmp31[179], tmp31[178], tmp31[177], tmp31[176], tmp31[175], tmp31[174], tmp31[173], tmp31[172], tmp31[171], tmp31[170], tmp31[169], tmp31[168], tmp31[167], tmp31[166], tmp31[165], tmp31[164], tmp31[163], tmp31[162], tmp31[161], tmp31[160], tmp31[159], tmp31[158], tmp31[157], tmp31[156], tmp31[155], tmp31[154], tmp31[153], tmp31[152], tmp31[151], tmp31[150], tmp31[149], tmp31[148], tmp31[147], tmp31[146], tmp31[145], tmp31[144], tmp31[143], tmp31[142], tmp31[141], tmp31[140], tmp31[139], tmp31[138], tmp31[137], tmp31[136], tmp31[135], tmp31[134], tmp31[133], tmp31[132], tmp31[131], tmp31[130], tmp31[129], tmp31[128], tmp31[127], tmp31[126], tmp31[125], tmp31[124], tmp31[123], tmp31[122], tmp31[121], tmp31[120], tmp31[119], tmp31[118], tmp31[117], tmp31[116], tmp31[115], tmp31[114], tmp31[113], tmp31[112], tmp31[111], tmp31[110], tmp31[109], tmp31[108], tmp31[107], tmp31[106], tmp31[105], tmp31[104], tmp31[103], tmp31[102], tmp31[101], tmp31[100], tmp31[99], tmp31[98], tmp31[97], tmp31[96], tmp31[95], tmp31[94], tmp31[93], tmp31[92], tmp31[91], tmp31[90], tmp31[89], tmp31[88], tmp31[87], tmp31[86], tmp31[85], tmp31[84], tmp31[83], tmp31[82], tmp31[81], tmp31[80], tmp31[79], tmp31[78], tmp31[77], tmp31[76], tmp31[75], tmp31[74], tmp31[73], tmp31[72], tmp31[71], tmp31[70], tmp31[69], tmp31[68], tmp31[67], tmp31[66], tmp31[65], tmp31[64], tmp31[63], tmp31[62], tmp31[61], tmp31[60], tmp31[59], tmp31[58], tmp31[57], tmp31[56], tmp31[55], tmp31[54], tmp31[53], tmp31[52], tmp31[51], tmp31[50], tmp31[49], tmp31[48], tmp31[47], tmp31[46], tmp31[45], tmp31[44], tmp31[43], tmp31[42], tmp31[41], tmp31[40], tmp31[39], tmp31[38], tmp31[37], tmp31[36], tmp31[35], tmp31[34], tmp31[33], tmp31[32], tmp31[31], tmp31[30], tmp31[29], tmp31[28], tmp31[27], tmp31[26], tmp31[25], tmp31[24], tmp31[23], tmp31[22], tmp31[21], tmp31[20], tmp31[19], tmp31[18], tmp31[17], tmp31[16], tmp31[15], tmp31[14], tmp31[13], tmp31[12], tmp31[11], tmp31[10], tmp31[9], tmp31[8], tmp31[7], tmp31[6], tmp31[5], tmp31[4], tmp31[3], tmp31[2], tmp31[1], tmp31[0]};
    assign tmp4368 = {tmp4367, const_417_0};
    assign tmp4369 = {const_418_0};
    assign tmp4370 = {tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369, tmp4369};
    assign tmp4371 = {tmp4370, const_418_0};
    assign tmp4372 = {tmp31[255]};
    assign tmp4373 = tmp4371 - tmp31;
    assign tmp4374 = {tmp4373[256]};
    assign tmp4375 = {tmp4371[255]};
    assign tmp4376 = ~tmp4375;
    assign tmp4377 = tmp4374 ^ tmp4376;
    assign tmp4378 = {tmp31[255]};
    assign tmp4379 = ~tmp4378;
    assign tmp4380 = tmp4377 ^ tmp4379;
    assign tmp4381 = {tmp4368[255]};
    assign tmp4382 = {const_419_0};
    assign tmp4383 = {tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382, tmp4382};
    assign tmp4384 = {tmp4383, const_419_0};
    assign tmp4385 = tmp4368 - tmp4384;
    assign tmp4386 = {tmp4385[256]};
    assign tmp4387 = {tmp4368[255]};
    assign tmp4388 = ~tmp4387;
    assign tmp4389 = tmp4386 ^ tmp4388;
    assign tmp4390 = {tmp4384[255]};
    assign tmp4391 = ~tmp4390;
    assign tmp4392 = tmp4389 ^ tmp4391;
    assign tmp4393 = tmp4380 & tmp4392;
    assign tmp4394 = {tmp31[255]};
    assign tmp4395 = {const_420_0};
    assign tmp4396 = {tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395, tmp4395};
    assign tmp4397 = {tmp4396, const_420_0};
    assign tmp4398 = tmp31 - tmp4397;
    assign tmp4399 = {tmp4398[256]};
    assign tmp4400 = {tmp31[255]};
    assign tmp4401 = ~tmp4400;
    assign tmp4402 = tmp4399 ^ tmp4401;
    assign tmp4403 = {tmp4397[255]};
    assign tmp4404 = ~tmp4403;
    assign tmp4405 = tmp4402 ^ tmp4404;
    assign tmp4406 = {const_421_0};
    assign tmp4407 = {tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406, tmp4406};
    assign tmp4408 = {tmp4407, const_421_0};
    assign tmp4409 = {tmp4368[255]};
    assign tmp4410 = tmp4408 - tmp4368;
    assign tmp4411 = {tmp4410[256]};
    assign tmp4412 = {tmp4408[255]};
    assign tmp4413 = ~tmp4412;
    assign tmp4414 = tmp4411 ^ tmp4413;
    assign tmp4415 = {tmp4368[255]};
    assign tmp4416 = ~tmp4415;
    assign tmp4417 = tmp4414 ^ tmp4416;
    assign tmp4418 = tmp4408 == tmp4368;
    assign tmp4419 = tmp4417 | tmp4418;
    assign tmp4420 = tmp4405 & tmp4419;
    assign tmp4421 = tmp4393 ? const_422_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp4368;
    assign tmp4422 = tmp4420 ? _ver_out_tmp_2 : tmp4421;
    assign tmp4423 = {tmp27[255]};
    assign tmp4424 = {tmp4422[255]};
    assign tmp4425 = tmp27 - tmp4422;
    assign tmp4426 = {tmp4425[256]};
    assign tmp4427 = {tmp27[255]};
    assign tmp4428 = ~tmp4427;
    assign tmp4429 = tmp4426 ^ tmp4428;
    assign tmp4430 = {tmp4422[255]};
    assign tmp4431 = ~tmp4430;
    assign tmp4432 = tmp4429 ^ tmp4431;
    assign tmp4433 = tmp4366 & tmp4432;
    assign tmp4434 = {tmp32[255]};
    assign tmp4435 = {tmp28[255]};
    assign tmp4436 = tmp32 - tmp28;
    assign tmp4437 = {tmp4436[256]};
    assign tmp4438 = {tmp32[255]};
    assign tmp4439 = ~tmp4438;
    assign tmp4440 = tmp4437 ^ tmp4439;
    assign tmp4441 = {tmp28[255]};
    assign tmp4442 = ~tmp4441;
    assign tmp4443 = tmp4440 ^ tmp4442;
    assign tmp4444 = tmp4433 & tmp4443;
    assign tmp4445 = {tmp32[253], tmp32[252], tmp32[251], tmp32[250], tmp32[249], tmp32[248], tmp32[247], tmp32[246], tmp32[245], tmp32[244], tmp32[243], tmp32[242], tmp32[241], tmp32[240], tmp32[239], tmp32[238], tmp32[237], tmp32[236], tmp32[235], tmp32[234], tmp32[233], tmp32[232], tmp32[231], tmp32[230], tmp32[229], tmp32[228], tmp32[227], tmp32[226], tmp32[225], tmp32[224], tmp32[223], tmp32[222], tmp32[221], tmp32[220], tmp32[219], tmp32[218], tmp32[217], tmp32[216], tmp32[215], tmp32[214], tmp32[213], tmp32[212], tmp32[211], tmp32[210], tmp32[209], tmp32[208], tmp32[207], tmp32[206], tmp32[205], tmp32[204], tmp32[203], tmp32[202], tmp32[201], tmp32[200], tmp32[199], tmp32[198], tmp32[197], tmp32[196], tmp32[195], tmp32[194], tmp32[193], tmp32[192], tmp32[191], tmp32[190], tmp32[189], tmp32[188], tmp32[187], tmp32[186], tmp32[185], tmp32[184], tmp32[183], tmp32[182], tmp32[181], tmp32[180], tmp32[179], tmp32[178], tmp32[177], tmp32[176], tmp32[175], tmp32[174], tmp32[173], tmp32[172], tmp32[171], tmp32[170], tmp32[169], tmp32[168], tmp32[167], tmp32[166], tmp32[165], tmp32[164], tmp32[163], tmp32[162], tmp32[161], tmp32[160], tmp32[159], tmp32[158], tmp32[157], tmp32[156], tmp32[155], tmp32[154], tmp32[153], tmp32[152], tmp32[151], tmp32[150], tmp32[149], tmp32[148], tmp32[147], tmp32[146], tmp32[145], tmp32[144], tmp32[143], tmp32[142], tmp32[141], tmp32[140], tmp32[139], tmp32[138], tmp32[137], tmp32[136], tmp32[135], tmp32[134], tmp32[133], tmp32[132], tmp32[131], tmp32[130], tmp32[129], tmp32[128], tmp32[127], tmp32[126], tmp32[125], tmp32[124], tmp32[123], tmp32[122], tmp32[121], tmp32[120], tmp32[119], tmp32[118], tmp32[117], tmp32[116], tmp32[115], tmp32[114], tmp32[113], tmp32[112], tmp32[111], tmp32[110], tmp32[109], tmp32[108], tmp32[107], tmp32[106], tmp32[105], tmp32[104], tmp32[103], tmp32[102], tmp32[101], tmp32[100], tmp32[99], tmp32[98], tmp32[97], tmp32[96], tmp32[95], tmp32[94], tmp32[93], tmp32[92], tmp32[91], tmp32[90], tmp32[89], tmp32[88], tmp32[87], tmp32[86], tmp32[85], tmp32[84], tmp32[83], tmp32[82], tmp32[81], tmp32[80], tmp32[79], tmp32[78], tmp32[77], tmp32[76], tmp32[75], tmp32[74], tmp32[73], tmp32[72], tmp32[71], tmp32[70], tmp32[69], tmp32[68], tmp32[67], tmp32[66], tmp32[65], tmp32[64], tmp32[63], tmp32[62], tmp32[61], tmp32[60], tmp32[59], tmp32[58], tmp32[57], tmp32[56], tmp32[55], tmp32[54], tmp32[53], tmp32[52], tmp32[51], tmp32[50], tmp32[49], tmp32[48], tmp32[47], tmp32[46], tmp32[45], tmp32[44], tmp32[43], tmp32[42], tmp32[41], tmp32[40], tmp32[39], tmp32[38], tmp32[37], tmp32[36], tmp32[35], tmp32[34], tmp32[33], tmp32[32], tmp32[31], tmp32[30], tmp32[29], tmp32[28], tmp32[27], tmp32[26], tmp32[25], tmp32[24], tmp32[23], tmp32[22], tmp32[21], tmp32[20], tmp32[19], tmp32[18], tmp32[17], tmp32[16], tmp32[15], tmp32[14], tmp32[13], tmp32[12], tmp32[11], tmp32[10], tmp32[9], tmp32[8], tmp32[7], tmp32[6], tmp32[5], tmp32[4], tmp32[3], tmp32[2], tmp32[1], tmp32[0]};
    assign tmp4446 = {tmp4445, const_424_0};
    assign tmp4447 = {const_425_0};
    assign tmp4448 = {tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447, tmp4447};
    assign tmp4449 = {tmp4448, const_425_0};
    assign tmp4450 = {tmp32[255]};
    assign tmp4451 = tmp4449 - tmp32;
    assign tmp4452 = {tmp4451[256]};
    assign tmp4453 = {tmp4449[255]};
    assign tmp4454 = ~tmp4453;
    assign tmp4455 = tmp4452 ^ tmp4454;
    assign tmp4456 = {tmp32[255]};
    assign tmp4457 = ~tmp4456;
    assign tmp4458 = tmp4455 ^ tmp4457;
    assign tmp4459 = {tmp4446[255]};
    assign tmp4460 = {const_426_0};
    assign tmp4461 = {tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460, tmp4460};
    assign tmp4462 = {tmp4461, const_426_0};
    assign tmp4463 = tmp4446 - tmp4462;
    assign tmp4464 = {tmp4463[256]};
    assign tmp4465 = {tmp4446[255]};
    assign tmp4466 = ~tmp4465;
    assign tmp4467 = tmp4464 ^ tmp4466;
    assign tmp4468 = {tmp4462[255]};
    assign tmp4469 = ~tmp4468;
    assign tmp4470 = tmp4467 ^ tmp4469;
    assign tmp4471 = tmp4458 & tmp4470;
    assign tmp4472 = {tmp32[255]};
    assign tmp4473 = {const_427_0};
    assign tmp4474 = {tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473, tmp4473};
    assign tmp4475 = {tmp4474, const_427_0};
    assign tmp4476 = tmp32 - tmp4475;
    assign tmp4477 = {tmp4476[256]};
    assign tmp4478 = {tmp32[255]};
    assign tmp4479 = ~tmp4478;
    assign tmp4480 = tmp4477 ^ tmp4479;
    assign tmp4481 = {tmp4475[255]};
    assign tmp4482 = ~tmp4481;
    assign tmp4483 = tmp4480 ^ tmp4482;
    assign tmp4484 = {const_428_0};
    assign tmp4485 = {tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484, tmp4484};
    assign tmp4486 = {tmp4485, const_428_0};
    assign tmp4487 = {tmp4446[255]};
    assign tmp4488 = tmp4486 - tmp4446;
    assign tmp4489 = {tmp4488[256]};
    assign tmp4490 = {tmp4486[255]};
    assign tmp4491 = ~tmp4490;
    assign tmp4492 = tmp4489 ^ tmp4491;
    assign tmp4493 = {tmp4446[255]};
    assign tmp4494 = ~tmp4493;
    assign tmp4495 = tmp4492 ^ tmp4494;
    assign tmp4496 = tmp4486 == tmp4446;
    assign tmp4497 = tmp4495 | tmp4496;
    assign tmp4498 = tmp4483 & tmp4497;
    assign tmp4499 = tmp4471 ? const_429_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp4446;
    assign tmp4500 = tmp4498 ? _ver_out_tmp_4 : tmp4499;
    assign tmp4501 = {tmp28[255]};
    assign tmp4502 = {tmp4500[255]};
    assign tmp4503 = tmp28 - tmp4500;
    assign tmp4504 = {tmp4503[256]};
    assign tmp4505 = {tmp28[255]};
    assign tmp4506 = ~tmp4505;
    assign tmp4507 = tmp4504 ^ tmp4506;
    assign tmp4508 = {tmp4500[255]};
    assign tmp4509 = ~tmp4508;
    assign tmp4510 = tmp4507 ^ tmp4509;
    assign tmp4511 = tmp4444 & tmp4510;
    assign tmp4512 = ~tmp35;
    assign tmp4513 = ~tmp36;
    assign tmp4514 = tmp4512 & tmp4513;
    assign tmp4515 = ~tmp57;
    assign tmp4516 = tmp4514 & tmp4515;
    assign tmp4517 = ~tmp1034;
    assign tmp4518 = tmp4516 & tmp4517;
    assign tmp4519 = tmp4518 & tmp2071;
    assign tmp4520 = ~tmp2583;
    assign tmp4521 = tmp4519 & tmp4520;
    assign tmp4522 = tmp4521 & tmp23;
    assign tmp4523 = ~tmp2627;
    assign tmp4524 = tmp4522 & tmp4523;
    assign tmp4525 = ~tmp2798;
    assign tmp4526 = tmp4524 & tmp4525;
    assign tmp4527 = ~tmp3425;
    assign tmp4528 = tmp4526 & tmp4527;
    assign tmp4529 = ~tmp4020;
    assign tmp4530 = tmp4528 & tmp4529;
    assign tmp4531 = tmp4530 & cfg_speculative_egest;
    assign tmp4532 = tmp4531 & tmp4511;
    assign tmp4533 = ~tmp35;
    assign tmp4534 = ~tmp36;
    assign tmp4535 = tmp4533 & tmp4534;
    assign tmp4536 = ~tmp57;
    assign tmp4537 = tmp4535 & tmp4536;
    assign tmp4538 = ~tmp1034;
    assign tmp4539 = tmp4537 & tmp4538;
    assign tmp4540 = tmp4539 & tmp2071;
    assign tmp4541 = ~tmp2583;
    assign tmp4542 = tmp4540 & tmp4541;
    assign tmp4543 = tmp4542 & tmp23;
    assign tmp4544 = ~tmp2627;
    assign tmp4545 = tmp4543 & tmp4544;
    assign tmp4546 = ~tmp2798;
    assign tmp4547 = tmp4545 & tmp4546;
    assign tmp4548 = ~tmp3425;
    assign tmp4549 = tmp4547 & tmp4548;
    assign tmp4550 = ~tmp4020;
    assign tmp4551 = tmp4549 & tmp4550;
    assign tmp4552 = tmp4551 & cfg_speculative_egest;
    assign tmp4553 = tmp4552 & tmp4511;
    assign tmp4554 = {tmp25[255], tmp25[254], tmp25[253], tmp25[252], tmp25[251], tmp25[250], tmp25[249], tmp25[248], tmp25[247], tmp25[246], tmp25[245], tmp25[244], tmp25[243], tmp25[242], tmp25[241], tmp25[240], tmp25[239], tmp25[238], tmp25[237], tmp25[236], tmp25[235], tmp25[234], tmp25[233], tmp25[232], tmp25[231], tmp25[230], tmp25[229], tmp25[228], tmp25[227], tmp25[226], tmp25[225], tmp25[224], tmp25[223], tmp25[222], tmp25[221], tmp25[220], tmp25[219], tmp25[218], tmp25[217], tmp25[216], tmp25[215], tmp25[214], tmp25[213], tmp25[212], tmp25[211], tmp25[210], tmp25[209], tmp25[208], tmp25[207], tmp25[206], tmp25[205], tmp25[204], tmp25[203], tmp25[202], tmp25[201], tmp25[200], tmp25[199], tmp25[198], tmp25[197], tmp25[196], tmp25[195], tmp25[194], tmp25[193], tmp25[192], tmp25[191], tmp25[190], tmp25[189], tmp25[188], tmp25[187], tmp25[186], tmp25[185], tmp25[184], tmp25[183], tmp25[182], tmp25[181], tmp25[180], tmp25[179], tmp25[178], tmp25[177], tmp25[176], tmp25[175], tmp25[174], tmp25[173], tmp25[172], tmp25[171], tmp25[170], tmp25[169], tmp25[168], tmp25[167], tmp25[166], tmp25[165], tmp25[164], tmp25[163], tmp25[162], tmp25[161], tmp25[160], tmp25[159], tmp25[158], tmp25[157], tmp25[156], tmp25[155], tmp25[154], tmp25[153], tmp25[152], tmp25[151], tmp25[150], tmp25[149], tmp25[148], tmp25[147], tmp25[146], tmp25[145], tmp25[144], tmp25[143], tmp25[142], tmp25[141], tmp25[140], tmp25[139], tmp25[138], tmp25[137], tmp25[136], tmp25[135], tmp25[134], tmp25[133], tmp25[132], tmp25[131], tmp25[130], tmp25[129], tmp25[128], tmp25[127], tmp25[126], tmp25[125], tmp25[124], tmp25[123], tmp25[122], tmp25[121], tmp25[120], tmp25[119], tmp25[118], tmp25[117], tmp25[116], tmp25[115], tmp25[114], tmp25[113], tmp25[112], tmp25[111], tmp25[110], tmp25[109], tmp25[108], tmp25[107], tmp25[106], tmp25[105], tmp25[104], tmp25[103], tmp25[102], tmp25[101], tmp25[100], tmp25[99], tmp25[98], tmp25[97], tmp25[96], tmp25[95], tmp25[94], tmp25[93], tmp25[92], tmp25[91], tmp25[90], tmp25[89], tmp25[88], tmp25[87], tmp25[86], tmp25[85], tmp25[84], tmp25[83], tmp25[82], tmp25[81], tmp25[80], tmp25[79], tmp25[78], tmp25[77], tmp25[76], tmp25[75], tmp25[74], tmp25[73], tmp25[72], tmp25[71], tmp25[70], tmp25[69], tmp25[68], tmp25[67], tmp25[66], tmp25[65], tmp25[64], tmp25[63], tmp25[62], tmp25[61], tmp25[60], tmp25[59], tmp25[58], tmp25[57], tmp25[56], tmp25[55], tmp25[54], tmp25[53], tmp25[52], tmp25[51], tmp25[50], tmp25[49], tmp25[48], tmp25[47], tmp25[46], tmp25[45], tmp25[44], tmp25[43], tmp25[42], tmp25[41], tmp25[40], tmp25[39], tmp25[38], tmp25[37], tmp25[36], tmp25[35], tmp25[34], tmp25[33], tmp25[32], tmp25[31], tmp25[30], tmp25[29], tmp25[28], tmp25[27], tmp25[26], tmp25[25], tmp25[24], tmp25[23], tmp25[22], tmp25[21], tmp25[20], tmp25[19], tmp25[18], tmp25[17], tmp25[16], tmp25[15], tmp25[14], tmp25[13], tmp25[12], tmp25[11], tmp25[10], tmp25[9], tmp25[8], tmp25[7], tmp25[6], tmp25[5], tmp25[4], tmp25[3], tmp25[2], tmp25[1]};
    assign tmp4555 = {tmp4554[254]};
    assign tmp4556 = {tmp4555};
    assign tmp4557 = {tmp4556, tmp4554};
    assign tmp4558 = ~tmp35;
    assign tmp4559 = ~tmp36;
    assign tmp4560 = tmp4558 & tmp4559;
    assign tmp4561 = ~tmp57;
    assign tmp4562 = tmp4560 & tmp4561;
    assign tmp4563 = ~tmp1034;
    assign tmp4564 = tmp4562 & tmp4563;
    assign tmp4565 = tmp4564 & tmp2071;
    assign tmp4566 = ~tmp2583;
    assign tmp4567 = tmp4565 & tmp4566;
    assign tmp4568 = tmp4567 & tmp23;
    assign tmp4569 = ~tmp2627;
    assign tmp4570 = tmp4568 & tmp4569;
    assign tmp4571 = ~tmp2798;
    assign tmp4572 = tmp4570 & tmp4571;
    assign tmp4573 = ~tmp3425;
    assign tmp4574 = tmp4572 & tmp4573;
    assign tmp4575 = ~tmp4020;
    assign tmp4576 = tmp4574 & tmp4575;
    assign tmp4577 = tmp4576 & cfg_speculative_egest;
    assign tmp4578 = tmp4577 & tmp4511;
    assign tmp4579 = tmp4578 & tmp24;
    assign tmp4580 = {tmp26[255], tmp26[254], tmp26[253], tmp26[252], tmp26[251], tmp26[250], tmp26[249], tmp26[248], tmp26[247], tmp26[246], tmp26[245], tmp26[244], tmp26[243], tmp26[242], tmp26[241], tmp26[240], tmp26[239], tmp26[238], tmp26[237], tmp26[236], tmp26[235], tmp26[234], tmp26[233], tmp26[232], tmp26[231], tmp26[230], tmp26[229], tmp26[228], tmp26[227], tmp26[226], tmp26[225], tmp26[224], tmp26[223], tmp26[222], tmp26[221], tmp26[220], tmp26[219], tmp26[218], tmp26[217], tmp26[216], tmp26[215], tmp26[214], tmp26[213], tmp26[212], tmp26[211], tmp26[210], tmp26[209], tmp26[208], tmp26[207], tmp26[206], tmp26[205], tmp26[204], tmp26[203], tmp26[202], tmp26[201], tmp26[200], tmp26[199], tmp26[198], tmp26[197], tmp26[196], tmp26[195], tmp26[194], tmp26[193], tmp26[192], tmp26[191], tmp26[190], tmp26[189], tmp26[188], tmp26[187], tmp26[186], tmp26[185], tmp26[184], tmp26[183], tmp26[182], tmp26[181], tmp26[180], tmp26[179], tmp26[178], tmp26[177], tmp26[176], tmp26[175], tmp26[174], tmp26[173], tmp26[172], tmp26[171], tmp26[170], tmp26[169], tmp26[168], tmp26[167], tmp26[166], tmp26[165], tmp26[164], tmp26[163], tmp26[162], tmp26[161], tmp26[160], tmp26[159], tmp26[158], tmp26[157], tmp26[156], tmp26[155], tmp26[154], tmp26[153], tmp26[152], tmp26[151], tmp26[150], tmp26[149], tmp26[148], tmp26[147], tmp26[146], tmp26[145], tmp26[144], tmp26[143], tmp26[142], tmp26[141], tmp26[140], tmp26[139], tmp26[138], tmp26[137], tmp26[136], tmp26[135], tmp26[134], tmp26[133], tmp26[132], tmp26[131], tmp26[130], tmp26[129], tmp26[128], tmp26[127], tmp26[126], tmp26[125], tmp26[124], tmp26[123], tmp26[122], tmp26[121], tmp26[120], tmp26[119], tmp26[118], tmp26[117], tmp26[116], tmp26[115], tmp26[114], tmp26[113], tmp26[112], tmp26[111], tmp26[110], tmp26[109], tmp26[108], tmp26[107], tmp26[106], tmp26[105], tmp26[104], tmp26[103], tmp26[102], tmp26[101], tmp26[100], tmp26[99], tmp26[98], tmp26[97], tmp26[96], tmp26[95], tmp26[94], tmp26[93], tmp26[92], tmp26[91], tmp26[90], tmp26[89], tmp26[88], tmp26[87], tmp26[86], tmp26[85], tmp26[84], tmp26[83], tmp26[82], tmp26[81], tmp26[80], tmp26[79], tmp26[78], tmp26[77], tmp26[76], tmp26[75], tmp26[74], tmp26[73], tmp26[72], tmp26[71], tmp26[70], tmp26[69], tmp26[68], tmp26[67], tmp26[66], tmp26[65], tmp26[64], tmp26[63], tmp26[62], tmp26[61], tmp26[60], tmp26[59], tmp26[58], tmp26[57], tmp26[56], tmp26[55], tmp26[54], tmp26[53], tmp26[52], tmp26[51], tmp26[50], tmp26[49], tmp26[48], tmp26[47], tmp26[46], tmp26[45], tmp26[44], tmp26[43], tmp26[42], tmp26[41], tmp26[40], tmp26[39], tmp26[38], tmp26[37], tmp26[36], tmp26[35], tmp26[34], tmp26[33], tmp26[32], tmp26[31], tmp26[30], tmp26[29], tmp26[28], tmp26[27], tmp26[26], tmp26[25], tmp26[24], tmp26[23], tmp26[22], tmp26[21], tmp26[20], tmp26[19], tmp26[18], tmp26[17], tmp26[16], tmp26[15], tmp26[14], tmp26[13], tmp26[12], tmp26[11], tmp26[10], tmp26[9], tmp26[8], tmp26[7], tmp26[6], tmp26[5], tmp26[4], tmp26[3], tmp26[2], tmp26[1]};
    assign tmp4581 = {tmp4580[254]};
    assign tmp4582 = {tmp4581};
    assign tmp4583 = {tmp4582, tmp4580};
    assign tmp4584 = ~tmp35;
    assign tmp4585 = ~tmp36;
    assign tmp4586 = tmp4584 & tmp4585;
    assign tmp4587 = ~tmp57;
    assign tmp4588 = tmp4586 & tmp4587;
    assign tmp4589 = ~tmp1034;
    assign tmp4590 = tmp4588 & tmp4589;
    assign tmp4591 = tmp4590 & tmp2071;
    assign tmp4592 = ~tmp2583;
    assign tmp4593 = tmp4591 & tmp4592;
    assign tmp4594 = tmp4593 & tmp23;
    assign tmp4595 = ~tmp2627;
    assign tmp4596 = tmp4594 & tmp4595;
    assign tmp4597 = ~tmp2798;
    assign tmp4598 = tmp4596 & tmp4597;
    assign tmp4599 = ~tmp3425;
    assign tmp4600 = tmp4598 & tmp4599;
    assign tmp4601 = ~tmp4020;
    assign tmp4602 = tmp4600 & tmp4601;
    assign tmp4603 = tmp4602 & cfg_speculative_egest;
    assign tmp4604 = tmp4603 & tmp4511;
    assign tmp4605 = tmp4604 & tmp24;
    assign tmp4606 = {tmp27[255], tmp27[254], tmp27[253], tmp27[252], tmp27[251], tmp27[250], tmp27[249], tmp27[248], tmp27[247], tmp27[246], tmp27[245], tmp27[244], tmp27[243], tmp27[242], tmp27[241], tmp27[240], tmp27[239], tmp27[238], tmp27[237], tmp27[236], tmp27[235], tmp27[234], tmp27[233], tmp27[232], tmp27[231], tmp27[230], tmp27[229], tmp27[228], tmp27[227], tmp27[226], tmp27[225], tmp27[224], tmp27[223], tmp27[222], tmp27[221], tmp27[220], tmp27[219], tmp27[218], tmp27[217], tmp27[216], tmp27[215], tmp27[214], tmp27[213], tmp27[212], tmp27[211], tmp27[210], tmp27[209], tmp27[208], tmp27[207], tmp27[206], tmp27[205], tmp27[204], tmp27[203], tmp27[202], tmp27[201], tmp27[200], tmp27[199], tmp27[198], tmp27[197], tmp27[196], tmp27[195], tmp27[194], tmp27[193], tmp27[192], tmp27[191], tmp27[190], tmp27[189], tmp27[188], tmp27[187], tmp27[186], tmp27[185], tmp27[184], tmp27[183], tmp27[182], tmp27[181], tmp27[180], tmp27[179], tmp27[178], tmp27[177], tmp27[176], tmp27[175], tmp27[174], tmp27[173], tmp27[172], tmp27[171], tmp27[170], tmp27[169], tmp27[168], tmp27[167], tmp27[166], tmp27[165], tmp27[164], tmp27[163], tmp27[162], tmp27[161], tmp27[160], tmp27[159], tmp27[158], tmp27[157], tmp27[156], tmp27[155], tmp27[154], tmp27[153], tmp27[152], tmp27[151], tmp27[150], tmp27[149], tmp27[148], tmp27[147], tmp27[146], tmp27[145], tmp27[144], tmp27[143], tmp27[142], tmp27[141], tmp27[140], tmp27[139], tmp27[138], tmp27[137], tmp27[136], tmp27[135], tmp27[134], tmp27[133], tmp27[132], tmp27[131], tmp27[130], tmp27[129], tmp27[128], tmp27[127], tmp27[126], tmp27[125], tmp27[124], tmp27[123], tmp27[122], tmp27[121], tmp27[120], tmp27[119], tmp27[118], tmp27[117], tmp27[116], tmp27[115], tmp27[114], tmp27[113], tmp27[112], tmp27[111], tmp27[110], tmp27[109], tmp27[108], tmp27[107], tmp27[106], tmp27[105], tmp27[104], tmp27[103], tmp27[102], tmp27[101], tmp27[100], tmp27[99], tmp27[98], tmp27[97], tmp27[96], tmp27[95], tmp27[94], tmp27[93], tmp27[92], tmp27[91], tmp27[90], tmp27[89], tmp27[88], tmp27[87], tmp27[86], tmp27[85], tmp27[84], tmp27[83], tmp27[82], tmp27[81], tmp27[80], tmp27[79], tmp27[78], tmp27[77], tmp27[76], tmp27[75], tmp27[74], tmp27[73], tmp27[72], tmp27[71], tmp27[70], tmp27[69], tmp27[68], tmp27[67], tmp27[66], tmp27[65], tmp27[64], tmp27[63], tmp27[62], tmp27[61], tmp27[60], tmp27[59], tmp27[58], tmp27[57], tmp27[56], tmp27[55], tmp27[54], tmp27[53], tmp27[52], tmp27[51], tmp27[50], tmp27[49], tmp27[48], tmp27[47], tmp27[46], tmp27[45], tmp27[44], tmp27[43], tmp27[42], tmp27[41], tmp27[40], tmp27[39], tmp27[38], tmp27[37], tmp27[36], tmp27[35], tmp27[34], tmp27[33], tmp27[32], tmp27[31], tmp27[30], tmp27[29], tmp27[28], tmp27[27], tmp27[26], tmp27[25], tmp27[24], tmp27[23], tmp27[22], tmp27[21], tmp27[20], tmp27[19], tmp27[18], tmp27[17], tmp27[16], tmp27[15], tmp27[14], tmp27[13], tmp27[12], tmp27[11], tmp27[10], tmp27[9], tmp27[8], tmp27[7], tmp27[6], tmp27[5], tmp27[4], tmp27[3], tmp27[2], tmp27[1]};
    assign tmp4607 = {tmp4606[254]};
    assign tmp4608 = {tmp4607};
    assign tmp4609 = {tmp4608, tmp4606};
    assign tmp4610 = ~tmp35;
    assign tmp4611 = ~tmp36;
    assign tmp4612 = tmp4610 & tmp4611;
    assign tmp4613 = ~tmp57;
    assign tmp4614 = tmp4612 & tmp4613;
    assign tmp4615 = ~tmp1034;
    assign tmp4616 = tmp4614 & tmp4615;
    assign tmp4617 = tmp4616 & tmp2071;
    assign tmp4618 = ~tmp2583;
    assign tmp4619 = tmp4617 & tmp4618;
    assign tmp4620 = tmp4619 & tmp23;
    assign tmp4621 = ~tmp2627;
    assign tmp4622 = tmp4620 & tmp4621;
    assign tmp4623 = ~tmp2798;
    assign tmp4624 = tmp4622 & tmp4623;
    assign tmp4625 = ~tmp3425;
    assign tmp4626 = tmp4624 & tmp4625;
    assign tmp4627 = ~tmp4020;
    assign tmp4628 = tmp4626 & tmp4627;
    assign tmp4629 = tmp4628 & cfg_speculative_egest;
    assign tmp4630 = tmp4629 & tmp4511;
    assign tmp4631 = tmp4630 & tmp24;
    assign tmp4632 = {tmp28[255], tmp28[254], tmp28[253], tmp28[252], tmp28[251], tmp28[250], tmp28[249], tmp28[248], tmp28[247], tmp28[246], tmp28[245], tmp28[244], tmp28[243], tmp28[242], tmp28[241], tmp28[240], tmp28[239], tmp28[238], tmp28[237], tmp28[236], tmp28[235], tmp28[234], tmp28[233], tmp28[232], tmp28[231], tmp28[230], tmp28[229], tmp28[228], tmp28[227], tmp28[226], tmp28[225], tmp28[224], tmp28[223], tmp28[222], tmp28[221], tmp28[220], tmp28[219], tmp28[218], tmp28[217], tmp28[216], tmp28[215], tmp28[214], tmp28[213], tmp28[212], tmp28[211], tmp28[210], tmp28[209], tmp28[208], tmp28[207], tmp28[206], tmp28[205], tmp28[204], tmp28[203], tmp28[202], tmp28[201], tmp28[200], tmp28[199], tmp28[198], tmp28[197], tmp28[196], tmp28[195], tmp28[194], tmp28[193], tmp28[192], tmp28[191], tmp28[190], tmp28[189], tmp28[188], tmp28[187], tmp28[186], tmp28[185], tmp28[184], tmp28[183], tmp28[182], tmp28[181], tmp28[180], tmp28[179], tmp28[178], tmp28[177], tmp28[176], tmp28[175], tmp28[174], tmp28[173], tmp28[172], tmp28[171], tmp28[170], tmp28[169], tmp28[168], tmp28[167], tmp28[166], tmp28[165], tmp28[164], tmp28[163], tmp28[162], tmp28[161], tmp28[160], tmp28[159], tmp28[158], tmp28[157], tmp28[156], tmp28[155], tmp28[154], tmp28[153], tmp28[152], tmp28[151], tmp28[150], tmp28[149], tmp28[148], tmp28[147], tmp28[146], tmp28[145], tmp28[144], tmp28[143], tmp28[142], tmp28[141], tmp28[140], tmp28[139], tmp28[138], tmp28[137], tmp28[136], tmp28[135], tmp28[134], tmp28[133], tmp28[132], tmp28[131], tmp28[130], tmp28[129], tmp28[128], tmp28[127], tmp28[126], tmp28[125], tmp28[124], tmp28[123], tmp28[122], tmp28[121], tmp28[120], tmp28[119], tmp28[118], tmp28[117], tmp28[116], tmp28[115], tmp28[114], tmp28[113], tmp28[112], tmp28[111], tmp28[110], tmp28[109], tmp28[108], tmp28[107], tmp28[106], tmp28[105], tmp28[104], tmp28[103], tmp28[102], tmp28[101], tmp28[100], tmp28[99], tmp28[98], tmp28[97], tmp28[96], tmp28[95], tmp28[94], tmp28[93], tmp28[92], tmp28[91], tmp28[90], tmp28[89], tmp28[88], tmp28[87], tmp28[86], tmp28[85], tmp28[84], tmp28[83], tmp28[82], tmp28[81], tmp28[80], tmp28[79], tmp28[78], tmp28[77], tmp28[76], tmp28[75], tmp28[74], tmp28[73], tmp28[72], tmp28[71], tmp28[70], tmp28[69], tmp28[68], tmp28[67], tmp28[66], tmp28[65], tmp28[64], tmp28[63], tmp28[62], tmp28[61], tmp28[60], tmp28[59], tmp28[58], tmp28[57], tmp28[56], tmp28[55], tmp28[54], tmp28[53], tmp28[52], tmp28[51], tmp28[50], tmp28[49], tmp28[48], tmp28[47], tmp28[46], tmp28[45], tmp28[44], tmp28[43], tmp28[42], tmp28[41], tmp28[40], tmp28[39], tmp28[38], tmp28[37], tmp28[36], tmp28[35], tmp28[34], tmp28[33], tmp28[32], tmp28[31], tmp28[30], tmp28[29], tmp28[28], tmp28[27], tmp28[26], tmp28[25], tmp28[24], tmp28[23], tmp28[22], tmp28[21], tmp28[20], tmp28[19], tmp28[18], tmp28[17], tmp28[16], tmp28[15], tmp28[14], tmp28[13], tmp28[12], tmp28[11], tmp28[10], tmp28[9], tmp28[8], tmp28[7], tmp28[6], tmp28[5], tmp28[4], tmp28[3], tmp28[2], tmp28[1]};
    assign tmp4633 = {tmp4632[254]};
    assign tmp4634 = {tmp4633};
    assign tmp4635 = {tmp4634, tmp4632};
    assign tmp4636 = ~tmp35;
    assign tmp4637 = ~tmp36;
    assign tmp4638 = tmp4636 & tmp4637;
    assign tmp4639 = ~tmp57;
    assign tmp4640 = tmp4638 & tmp4639;
    assign tmp4641 = ~tmp1034;
    assign tmp4642 = tmp4640 & tmp4641;
    assign tmp4643 = tmp4642 & tmp2071;
    assign tmp4644 = ~tmp2583;
    assign tmp4645 = tmp4643 & tmp4644;
    assign tmp4646 = tmp4645 & tmp23;
    assign tmp4647 = ~tmp2627;
    assign tmp4648 = tmp4646 & tmp4647;
    assign tmp4649 = ~tmp2798;
    assign tmp4650 = tmp4648 & tmp4649;
    assign tmp4651 = ~tmp3425;
    assign tmp4652 = tmp4650 & tmp4651;
    assign tmp4653 = ~tmp4020;
    assign tmp4654 = tmp4652 & tmp4653;
    assign tmp4655 = tmp4654 & cfg_speculative_egest;
    assign tmp4656 = tmp4655 & tmp4511;
    assign tmp4657 = tmp4656 & tmp24;
    assign tmp4658 = ~tmp35;
    assign tmp4659 = ~tmp36;
    assign tmp4660 = tmp4658 & tmp4659;
    assign tmp4661 = ~tmp57;
    assign tmp4662 = tmp4660 & tmp4661;
    assign tmp4663 = ~tmp1034;
    assign tmp4664 = tmp4662 & tmp4663;
    assign tmp4665 = tmp4664 & tmp2071;
    assign tmp4666 = ~tmp2583;
    assign tmp4667 = tmp4665 & tmp4666;
    assign tmp4668 = tmp4667 & tmp23;
    assign tmp4669 = ~tmp2627;
    assign tmp4670 = tmp4668 & tmp4669;
    assign tmp4671 = ~tmp2798;
    assign tmp4672 = tmp4670 & tmp4671;
    assign tmp4673 = ~tmp3425;
    assign tmp4674 = tmp4672 & tmp4673;
    assign tmp4675 = ~tmp4020;
    assign tmp4676 = tmp4674 & tmp4675;
    assign tmp4677 = tmp4676 & cfg_speculative_egest;
    assign tmp4678 = tmp4677 & tmp4511;
    assign tmp4679 = tmp4678 & tmp24;
    assign tmp4680 = ~tmp35;
    assign tmp4681 = ~tmp36;
    assign tmp4682 = tmp4680 & tmp4681;
    assign tmp4683 = ~tmp57;
    assign tmp4684 = tmp4682 & tmp4683;
    assign tmp4685 = ~tmp1034;
    assign tmp4686 = tmp4684 & tmp4685;
    assign tmp4687 = tmp4686 & tmp2071;
    assign tmp4688 = ~tmp2583;
    assign tmp4689 = tmp4687 & tmp4688;
    assign tmp4690 = tmp4689 & tmp23;
    assign tmp4691 = ~tmp2627;
    assign tmp4692 = tmp4690 & tmp4691;
    assign tmp4693 = ~tmp2798;
    assign tmp4694 = tmp4692 & tmp4693;
    assign tmp4695 = ~tmp3425;
    assign tmp4696 = tmp4694 & tmp4695;
    assign tmp4697 = ~tmp4020;
    assign tmp4698 = tmp4696 & tmp4697;
    assign tmp4699 = tmp4698 & cfg_speculative_egest;
    assign tmp4700 = tmp4699 & tmp4511;
    assign tmp4701 = tmp4700 & tmp24;
    assign tmp4702 = ~tmp35;
    assign tmp4703 = ~tmp36;
    assign tmp4704 = tmp4702 & tmp4703;
    assign tmp4705 = ~tmp57;
    assign tmp4706 = tmp4704 & tmp4705;
    assign tmp4707 = ~tmp1034;
    assign tmp4708 = tmp4706 & tmp4707;
    assign tmp4709 = tmp4708 & tmp2071;
    assign tmp4710 = ~tmp2583;
    assign tmp4711 = tmp4709 & tmp4710;
    assign tmp4712 = tmp4711 & tmp23;
    assign tmp4713 = ~tmp2627;
    assign tmp4714 = tmp4712 & tmp4713;
    assign tmp4715 = ~tmp2798;
    assign tmp4716 = tmp4714 & tmp4715;
    assign tmp4717 = ~tmp3425;
    assign tmp4718 = tmp4716 & tmp4717;
    assign tmp4719 = ~tmp4020;
    assign tmp4720 = tmp4718 & tmp4719;
    assign tmp4721 = tmp4720 & cfg_speculative_egest;
    assign tmp4722 = tmp4721 & tmp4511;
    assign tmp4723 = tmp4722 & tmp24;
    assign tmp4724 = ~tmp35;
    assign tmp4725 = ~tmp36;
    assign tmp4726 = tmp4724 & tmp4725;
    assign tmp4727 = ~tmp57;
    assign tmp4728 = tmp4726 & tmp4727;
    assign tmp4729 = ~tmp1034;
    assign tmp4730 = tmp4728 & tmp4729;
    assign tmp4731 = tmp4730 & tmp2071;
    assign tmp4732 = ~tmp2583;
    assign tmp4733 = tmp4731 & tmp4732;
    assign tmp4734 = tmp4733 & tmp23;
    assign tmp4735 = ~tmp2627;
    assign tmp4736 = tmp4734 & tmp4735;
    assign tmp4737 = ~tmp2798;
    assign tmp4738 = tmp4736 & tmp4737;
    assign tmp4739 = ~tmp3425;
    assign tmp4740 = tmp4738 & tmp4739;
    assign tmp4741 = ~tmp4020;
    assign tmp4742 = tmp4740 & tmp4741;
    assign tmp4743 = tmp4742 & cfg_speculative_egest;
    assign tmp4744 = tmp4743 & tmp4511;
    assign tmp4745 = tmp4744 & tmp24;
    assign tmp4746 = ~tmp35;
    assign tmp4747 = ~tmp36;
    assign tmp4748 = tmp4746 & tmp4747;
    assign tmp4749 = ~tmp57;
    assign tmp4750 = tmp4748 & tmp4749;
    assign tmp4751 = ~tmp1034;
    assign tmp4752 = tmp4750 & tmp4751;
    assign tmp4753 = tmp4752 & tmp2071;
    assign tmp4754 = ~tmp2583;
    assign tmp4755 = tmp4753 & tmp4754;
    assign tmp4756 = tmp4755 & tmp23;
    assign tmp4757 = ~tmp2627;
    assign tmp4758 = tmp4756 & tmp4757;
    assign tmp4759 = ~tmp2798;
    assign tmp4760 = tmp4758 & tmp4759;
    assign tmp4761 = ~tmp3425;
    assign tmp4762 = tmp4760 & tmp4761;
    assign tmp4763 = ~tmp4020;
    assign tmp4764 = tmp4762 & tmp4763;
    assign tmp4765 = tmp4764 & cfg_speculative_egest;
    assign tmp4766 = tmp4765 & tmp4511;
    assign tmp4767 = ~tmp24;
    assign tmp4768 = tmp4766 & tmp4767;
    assign tmp4769 = ~tmp35;
    assign tmp4770 = ~tmp36;
    assign tmp4771 = tmp4769 & tmp4770;
    assign tmp4772 = ~tmp57;
    assign tmp4773 = tmp4771 & tmp4772;
    assign tmp4774 = ~tmp1034;
    assign tmp4775 = tmp4773 & tmp4774;
    assign tmp4776 = tmp4775 & tmp2071;
    assign tmp4777 = ~tmp2583;
    assign tmp4778 = tmp4776 & tmp4777;
    assign tmp4779 = tmp4778 & tmp23;
    assign tmp4780 = ~tmp2627;
    assign tmp4781 = tmp4779 & tmp4780;
    assign tmp4782 = ~tmp2798;
    assign tmp4783 = tmp4781 & tmp4782;
    assign tmp4784 = ~tmp3425;
    assign tmp4785 = tmp4783 & tmp4784;
    assign tmp4786 = ~tmp4020;
    assign tmp4787 = tmp4785 & tmp4786;
    assign tmp4788 = tmp4787 & cfg_speculative_egest;
    assign tmp4789 = tmp4788 & tmp4511;
    assign tmp4790 = ~tmp24;
    assign tmp4791 = tmp4789 & tmp4790;
    assign tmp4792 = ~tmp35;
    assign tmp4793 = ~tmp36;
    assign tmp4794 = tmp4792 & tmp4793;
    assign tmp4795 = ~tmp57;
    assign tmp4796 = tmp4794 & tmp4795;
    assign tmp4797 = ~tmp1034;
    assign tmp4798 = tmp4796 & tmp4797;
    assign tmp4799 = tmp4798 & tmp2071;
    assign tmp4800 = ~tmp2583;
    assign tmp4801 = tmp4799 & tmp4800;
    assign tmp4802 = tmp4801 & tmp23;
    assign tmp4803 = ~tmp2627;
    assign tmp4804 = tmp4802 & tmp4803;
    assign tmp4805 = ~tmp2798;
    assign tmp4806 = tmp4804 & tmp4805;
    assign tmp4807 = ~tmp3425;
    assign tmp4808 = tmp4806 & tmp4807;
    assign tmp4809 = ~tmp4020;
    assign tmp4810 = tmp4808 & tmp4809;
    assign tmp4811 = tmp4810 & cfg_speculative_egest;
    assign tmp4812 = tmp4811 & tmp4511;
    assign tmp4813 = ~tmp24;
    assign tmp4814 = tmp4812 & tmp4813;
    assign tmp4815 = ~tmp35;
    assign tmp4816 = ~tmp36;
    assign tmp4817 = tmp4815 & tmp4816;
    assign tmp4818 = ~tmp57;
    assign tmp4819 = tmp4817 & tmp4818;
    assign tmp4820 = ~tmp1034;
    assign tmp4821 = tmp4819 & tmp4820;
    assign tmp4822 = tmp4821 & tmp2071;
    assign tmp4823 = ~tmp2583;
    assign tmp4824 = tmp4822 & tmp4823;
    assign tmp4825 = tmp4824 & tmp23;
    assign tmp4826 = ~tmp2627;
    assign tmp4827 = tmp4825 & tmp4826;
    assign tmp4828 = ~tmp2798;
    assign tmp4829 = tmp4827 & tmp4828;
    assign tmp4830 = ~tmp3425;
    assign tmp4831 = tmp4829 & tmp4830;
    assign tmp4832 = ~tmp4020;
    assign tmp4833 = tmp4831 & tmp4832;
    assign tmp4834 = tmp4833 & cfg_speculative_egest;
    assign tmp4835 = tmp4834 & tmp4511;
    assign tmp4836 = ~tmp24;
    assign tmp4837 = tmp4835 & tmp4836;
    assign tmp4838 = {tmp29[254], tmp29[253], tmp29[252], tmp29[251], tmp29[250], tmp29[249], tmp29[248], tmp29[247], tmp29[246], tmp29[245], tmp29[244], tmp29[243], tmp29[242], tmp29[241], tmp29[240], tmp29[239], tmp29[238], tmp29[237], tmp29[236], tmp29[235], tmp29[234], tmp29[233], tmp29[232], tmp29[231], tmp29[230], tmp29[229], tmp29[228], tmp29[227], tmp29[226], tmp29[225], tmp29[224], tmp29[223], tmp29[222], tmp29[221], tmp29[220], tmp29[219], tmp29[218], tmp29[217], tmp29[216], tmp29[215], tmp29[214], tmp29[213], tmp29[212], tmp29[211], tmp29[210], tmp29[209], tmp29[208], tmp29[207], tmp29[206], tmp29[205], tmp29[204], tmp29[203], tmp29[202], tmp29[201], tmp29[200], tmp29[199], tmp29[198], tmp29[197], tmp29[196], tmp29[195], tmp29[194], tmp29[193], tmp29[192], tmp29[191], tmp29[190], tmp29[189], tmp29[188], tmp29[187], tmp29[186], tmp29[185], tmp29[184], tmp29[183], tmp29[182], tmp29[181], tmp29[180], tmp29[179], tmp29[178], tmp29[177], tmp29[176], tmp29[175], tmp29[174], tmp29[173], tmp29[172], tmp29[171], tmp29[170], tmp29[169], tmp29[168], tmp29[167], tmp29[166], tmp29[165], tmp29[164], tmp29[163], tmp29[162], tmp29[161], tmp29[160], tmp29[159], tmp29[158], tmp29[157], tmp29[156], tmp29[155], tmp29[154], tmp29[153], tmp29[152], tmp29[151], tmp29[150], tmp29[149], tmp29[148], tmp29[147], tmp29[146], tmp29[145], tmp29[144], tmp29[143], tmp29[142], tmp29[141], tmp29[140], tmp29[139], tmp29[138], tmp29[137], tmp29[136], tmp29[135], tmp29[134], tmp29[133], tmp29[132], tmp29[131], tmp29[130], tmp29[129], tmp29[128], tmp29[127], tmp29[126], tmp29[125], tmp29[124], tmp29[123], tmp29[122], tmp29[121], tmp29[120], tmp29[119], tmp29[118], tmp29[117], tmp29[116], tmp29[115], tmp29[114], tmp29[113], tmp29[112], tmp29[111], tmp29[110], tmp29[109], tmp29[108], tmp29[107], tmp29[106], tmp29[105], tmp29[104], tmp29[103], tmp29[102], tmp29[101], tmp29[100], tmp29[99], tmp29[98], tmp29[97], tmp29[96], tmp29[95], tmp29[94], tmp29[93], tmp29[92], tmp29[91], tmp29[90], tmp29[89], tmp29[88], tmp29[87], tmp29[86], tmp29[85], tmp29[84], tmp29[83], tmp29[82], tmp29[81], tmp29[80], tmp29[79], tmp29[78], tmp29[77], tmp29[76], tmp29[75], tmp29[74], tmp29[73], tmp29[72], tmp29[71], tmp29[70], tmp29[69], tmp29[68], tmp29[67], tmp29[66], tmp29[65], tmp29[64], tmp29[63], tmp29[62], tmp29[61], tmp29[60], tmp29[59], tmp29[58], tmp29[57], tmp29[56], tmp29[55], tmp29[54], tmp29[53], tmp29[52], tmp29[51], tmp29[50], tmp29[49], tmp29[48], tmp29[47], tmp29[46], tmp29[45], tmp29[44], tmp29[43], tmp29[42], tmp29[41], tmp29[40], tmp29[39], tmp29[38], tmp29[37], tmp29[36], tmp29[35], tmp29[34], tmp29[33], tmp29[32], tmp29[31], tmp29[30], tmp29[29], tmp29[28], tmp29[27], tmp29[26], tmp29[25], tmp29[24], tmp29[23], tmp29[22], tmp29[21], tmp29[20], tmp29[19], tmp29[18], tmp29[17], tmp29[16], tmp29[15], tmp29[14], tmp29[13], tmp29[12], tmp29[11], tmp29[10], tmp29[9], tmp29[8], tmp29[7], tmp29[6], tmp29[5], tmp29[4], tmp29[3], tmp29[2], tmp29[1], tmp29[0]};
    assign tmp4839 = {tmp4838, const_433_0};
    assign tmp4840 = {const_434_0};
    assign tmp4841 = {tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840, tmp4840};
    assign tmp4842 = {tmp4841, const_434_0};
    assign tmp4843 = {tmp29[255]};
    assign tmp4844 = tmp4842 - tmp29;
    assign tmp4845 = {tmp4844[256]};
    assign tmp4846 = {tmp4842[255]};
    assign tmp4847 = ~tmp4846;
    assign tmp4848 = tmp4845 ^ tmp4847;
    assign tmp4849 = {tmp29[255]};
    assign tmp4850 = ~tmp4849;
    assign tmp4851 = tmp4848 ^ tmp4850;
    assign tmp4852 = {tmp4839[255]};
    assign tmp4853 = {const_435_0};
    assign tmp4854 = {tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853, tmp4853};
    assign tmp4855 = {tmp4854, const_435_0};
    assign tmp4856 = tmp4839 - tmp4855;
    assign tmp4857 = {tmp4856[256]};
    assign tmp4858 = {tmp4839[255]};
    assign tmp4859 = ~tmp4858;
    assign tmp4860 = tmp4857 ^ tmp4859;
    assign tmp4861 = {tmp4855[255]};
    assign tmp4862 = ~tmp4861;
    assign tmp4863 = tmp4860 ^ tmp4862;
    assign tmp4864 = tmp4851 & tmp4863;
    assign tmp4865 = {tmp29[255]};
    assign tmp4866 = {const_436_0};
    assign tmp4867 = {tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866, tmp4866};
    assign tmp4868 = {tmp4867, const_436_0};
    assign tmp4869 = tmp29 - tmp4868;
    assign tmp4870 = {tmp4869[256]};
    assign tmp4871 = {tmp29[255]};
    assign tmp4872 = ~tmp4871;
    assign tmp4873 = tmp4870 ^ tmp4872;
    assign tmp4874 = {tmp4868[255]};
    assign tmp4875 = ~tmp4874;
    assign tmp4876 = tmp4873 ^ tmp4875;
    assign tmp4877 = {const_437_0};
    assign tmp4878 = {tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877, tmp4877};
    assign tmp4879 = {tmp4878, const_437_0};
    assign tmp4880 = {tmp4839[255]};
    assign tmp4881 = tmp4879 - tmp4839;
    assign tmp4882 = {tmp4881[256]};
    assign tmp4883 = {tmp4879[255]};
    assign tmp4884 = ~tmp4883;
    assign tmp4885 = tmp4882 ^ tmp4884;
    assign tmp4886 = {tmp4839[255]};
    assign tmp4887 = ~tmp4886;
    assign tmp4888 = tmp4885 ^ tmp4887;
    assign tmp4889 = tmp4879 == tmp4839;
    assign tmp4890 = tmp4888 | tmp4889;
    assign tmp4891 = tmp4876 & tmp4890;
    assign tmp4892 = tmp4864 ? const_438_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp4839;
    assign tmp4893 = tmp4891 ? _ver_out_tmp_7 : tmp4892;
    assign tmp4894 = ~tmp35;
    assign tmp4895 = ~tmp36;
    assign tmp4896 = tmp4894 & tmp4895;
    assign tmp4897 = ~tmp57;
    assign tmp4898 = tmp4896 & tmp4897;
    assign tmp4899 = ~tmp1034;
    assign tmp4900 = tmp4898 & tmp4899;
    assign tmp4901 = tmp4900 & tmp2071;
    assign tmp4902 = ~tmp2583;
    assign tmp4903 = tmp4901 & tmp4902;
    assign tmp4904 = tmp4903 & tmp23;
    assign tmp4905 = ~tmp2627;
    assign tmp4906 = tmp4904 & tmp4905;
    assign tmp4907 = ~tmp2798;
    assign tmp4908 = tmp4906 & tmp4907;
    assign tmp4909 = ~tmp3425;
    assign tmp4910 = tmp4908 & tmp4909;
    assign tmp4911 = ~tmp4020;
    assign tmp4912 = tmp4910 & tmp4911;
    assign tmp4913 = tmp4912 & cfg_speculative_egest;
    assign tmp4914 = tmp4913 & tmp4511;
    assign tmp4915 = ~tmp24;
    assign tmp4916 = tmp4914 & tmp4915;
    assign tmp4917 = {tmp30[254], tmp30[253], tmp30[252], tmp30[251], tmp30[250], tmp30[249], tmp30[248], tmp30[247], tmp30[246], tmp30[245], tmp30[244], tmp30[243], tmp30[242], tmp30[241], tmp30[240], tmp30[239], tmp30[238], tmp30[237], tmp30[236], tmp30[235], tmp30[234], tmp30[233], tmp30[232], tmp30[231], tmp30[230], tmp30[229], tmp30[228], tmp30[227], tmp30[226], tmp30[225], tmp30[224], tmp30[223], tmp30[222], tmp30[221], tmp30[220], tmp30[219], tmp30[218], tmp30[217], tmp30[216], tmp30[215], tmp30[214], tmp30[213], tmp30[212], tmp30[211], tmp30[210], tmp30[209], tmp30[208], tmp30[207], tmp30[206], tmp30[205], tmp30[204], tmp30[203], tmp30[202], tmp30[201], tmp30[200], tmp30[199], tmp30[198], tmp30[197], tmp30[196], tmp30[195], tmp30[194], tmp30[193], tmp30[192], tmp30[191], tmp30[190], tmp30[189], tmp30[188], tmp30[187], tmp30[186], tmp30[185], tmp30[184], tmp30[183], tmp30[182], tmp30[181], tmp30[180], tmp30[179], tmp30[178], tmp30[177], tmp30[176], tmp30[175], tmp30[174], tmp30[173], tmp30[172], tmp30[171], tmp30[170], tmp30[169], tmp30[168], tmp30[167], tmp30[166], tmp30[165], tmp30[164], tmp30[163], tmp30[162], tmp30[161], tmp30[160], tmp30[159], tmp30[158], tmp30[157], tmp30[156], tmp30[155], tmp30[154], tmp30[153], tmp30[152], tmp30[151], tmp30[150], tmp30[149], tmp30[148], tmp30[147], tmp30[146], tmp30[145], tmp30[144], tmp30[143], tmp30[142], tmp30[141], tmp30[140], tmp30[139], tmp30[138], tmp30[137], tmp30[136], tmp30[135], tmp30[134], tmp30[133], tmp30[132], tmp30[131], tmp30[130], tmp30[129], tmp30[128], tmp30[127], tmp30[126], tmp30[125], tmp30[124], tmp30[123], tmp30[122], tmp30[121], tmp30[120], tmp30[119], tmp30[118], tmp30[117], tmp30[116], tmp30[115], tmp30[114], tmp30[113], tmp30[112], tmp30[111], tmp30[110], tmp30[109], tmp30[108], tmp30[107], tmp30[106], tmp30[105], tmp30[104], tmp30[103], tmp30[102], tmp30[101], tmp30[100], tmp30[99], tmp30[98], tmp30[97], tmp30[96], tmp30[95], tmp30[94], tmp30[93], tmp30[92], tmp30[91], tmp30[90], tmp30[89], tmp30[88], tmp30[87], tmp30[86], tmp30[85], tmp30[84], tmp30[83], tmp30[82], tmp30[81], tmp30[80], tmp30[79], tmp30[78], tmp30[77], tmp30[76], tmp30[75], tmp30[74], tmp30[73], tmp30[72], tmp30[71], tmp30[70], tmp30[69], tmp30[68], tmp30[67], tmp30[66], tmp30[65], tmp30[64], tmp30[63], tmp30[62], tmp30[61], tmp30[60], tmp30[59], tmp30[58], tmp30[57], tmp30[56], tmp30[55], tmp30[54], tmp30[53], tmp30[52], tmp30[51], tmp30[50], tmp30[49], tmp30[48], tmp30[47], tmp30[46], tmp30[45], tmp30[44], tmp30[43], tmp30[42], tmp30[41], tmp30[40], tmp30[39], tmp30[38], tmp30[37], tmp30[36], tmp30[35], tmp30[34], tmp30[33], tmp30[32], tmp30[31], tmp30[30], tmp30[29], tmp30[28], tmp30[27], tmp30[26], tmp30[25], tmp30[24], tmp30[23], tmp30[22], tmp30[21], tmp30[20], tmp30[19], tmp30[18], tmp30[17], tmp30[16], tmp30[15], tmp30[14], tmp30[13], tmp30[12], tmp30[11], tmp30[10], tmp30[9], tmp30[8], tmp30[7], tmp30[6], tmp30[5], tmp30[4], tmp30[3], tmp30[2], tmp30[1], tmp30[0]};
    assign tmp4918 = {tmp4917, const_440_0};
    assign tmp4919 = {const_441_0};
    assign tmp4920 = {tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919, tmp4919};
    assign tmp4921 = {tmp4920, const_441_0};
    assign tmp4922 = {tmp30[255]};
    assign tmp4923 = tmp4921 - tmp30;
    assign tmp4924 = {tmp4923[256]};
    assign tmp4925 = {tmp4921[255]};
    assign tmp4926 = ~tmp4925;
    assign tmp4927 = tmp4924 ^ tmp4926;
    assign tmp4928 = {tmp30[255]};
    assign tmp4929 = ~tmp4928;
    assign tmp4930 = tmp4927 ^ tmp4929;
    assign tmp4931 = {tmp4918[255]};
    assign tmp4932 = {const_442_0};
    assign tmp4933 = {tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932, tmp4932};
    assign tmp4934 = {tmp4933, const_442_0};
    assign tmp4935 = tmp4918 - tmp4934;
    assign tmp4936 = {tmp4935[256]};
    assign tmp4937 = {tmp4918[255]};
    assign tmp4938 = ~tmp4937;
    assign tmp4939 = tmp4936 ^ tmp4938;
    assign tmp4940 = {tmp4934[255]};
    assign tmp4941 = ~tmp4940;
    assign tmp4942 = tmp4939 ^ tmp4941;
    assign tmp4943 = tmp4930 & tmp4942;
    assign tmp4944 = {tmp30[255]};
    assign tmp4945 = {const_443_0};
    assign tmp4946 = {tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945, tmp4945};
    assign tmp4947 = {tmp4946, const_443_0};
    assign tmp4948 = tmp30 - tmp4947;
    assign tmp4949 = {tmp4948[256]};
    assign tmp4950 = {tmp30[255]};
    assign tmp4951 = ~tmp4950;
    assign tmp4952 = tmp4949 ^ tmp4951;
    assign tmp4953 = {tmp4947[255]};
    assign tmp4954 = ~tmp4953;
    assign tmp4955 = tmp4952 ^ tmp4954;
    assign tmp4956 = {const_444_0};
    assign tmp4957 = {tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956, tmp4956};
    assign tmp4958 = {tmp4957, const_444_0};
    assign tmp4959 = {tmp4918[255]};
    assign tmp4960 = tmp4958 - tmp4918;
    assign tmp4961 = {tmp4960[256]};
    assign tmp4962 = {tmp4958[255]};
    assign tmp4963 = ~tmp4962;
    assign tmp4964 = tmp4961 ^ tmp4963;
    assign tmp4965 = {tmp4918[255]};
    assign tmp4966 = ~tmp4965;
    assign tmp4967 = tmp4964 ^ tmp4966;
    assign tmp4968 = tmp4958 == tmp4918;
    assign tmp4969 = tmp4967 | tmp4968;
    assign tmp4970 = tmp4955 & tmp4969;
    assign tmp4971 = tmp4943 ? const_445_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp4918;
    assign tmp4972 = tmp4970 ? _ver_out_tmp_9 : tmp4971;
    assign tmp4973 = ~tmp35;
    assign tmp4974 = ~tmp36;
    assign tmp4975 = tmp4973 & tmp4974;
    assign tmp4976 = ~tmp57;
    assign tmp4977 = tmp4975 & tmp4976;
    assign tmp4978 = ~tmp1034;
    assign tmp4979 = tmp4977 & tmp4978;
    assign tmp4980 = tmp4979 & tmp2071;
    assign tmp4981 = ~tmp2583;
    assign tmp4982 = tmp4980 & tmp4981;
    assign tmp4983 = tmp4982 & tmp23;
    assign tmp4984 = ~tmp2627;
    assign tmp4985 = tmp4983 & tmp4984;
    assign tmp4986 = ~tmp2798;
    assign tmp4987 = tmp4985 & tmp4986;
    assign tmp4988 = ~tmp3425;
    assign tmp4989 = tmp4987 & tmp4988;
    assign tmp4990 = ~tmp4020;
    assign tmp4991 = tmp4989 & tmp4990;
    assign tmp4992 = tmp4991 & cfg_speculative_egest;
    assign tmp4993 = tmp4992 & tmp4511;
    assign tmp4994 = ~tmp24;
    assign tmp4995 = tmp4993 & tmp4994;
    assign tmp4996 = {tmp31[254], tmp31[253], tmp31[252], tmp31[251], tmp31[250], tmp31[249], tmp31[248], tmp31[247], tmp31[246], tmp31[245], tmp31[244], tmp31[243], tmp31[242], tmp31[241], tmp31[240], tmp31[239], tmp31[238], tmp31[237], tmp31[236], tmp31[235], tmp31[234], tmp31[233], tmp31[232], tmp31[231], tmp31[230], tmp31[229], tmp31[228], tmp31[227], tmp31[226], tmp31[225], tmp31[224], tmp31[223], tmp31[222], tmp31[221], tmp31[220], tmp31[219], tmp31[218], tmp31[217], tmp31[216], tmp31[215], tmp31[214], tmp31[213], tmp31[212], tmp31[211], tmp31[210], tmp31[209], tmp31[208], tmp31[207], tmp31[206], tmp31[205], tmp31[204], tmp31[203], tmp31[202], tmp31[201], tmp31[200], tmp31[199], tmp31[198], tmp31[197], tmp31[196], tmp31[195], tmp31[194], tmp31[193], tmp31[192], tmp31[191], tmp31[190], tmp31[189], tmp31[188], tmp31[187], tmp31[186], tmp31[185], tmp31[184], tmp31[183], tmp31[182], tmp31[181], tmp31[180], tmp31[179], tmp31[178], tmp31[177], tmp31[176], tmp31[175], tmp31[174], tmp31[173], tmp31[172], tmp31[171], tmp31[170], tmp31[169], tmp31[168], tmp31[167], tmp31[166], tmp31[165], tmp31[164], tmp31[163], tmp31[162], tmp31[161], tmp31[160], tmp31[159], tmp31[158], tmp31[157], tmp31[156], tmp31[155], tmp31[154], tmp31[153], tmp31[152], tmp31[151], tmp31[150], tmp31[149], tmp31[148], tmp31[147], tmp31[146], tmp31[145], tmp31[144], tmp31[143], tmp31[142], tmp31[141], tmp31[140], tmp31[139], tmp31[138], tmp31[137], tmp31[136], tmp31[135], tmp31[134], tmp31[133], tmp31[132], tmp31[131], tmp31[130], tmp31[129], tmp31[128], tmp31[127], tmp31[126], tmp31[125], tmp31[124], tmp31[123], tmp31[122], tmp31[121], tmp31[120], tmp31[119], tmp31[118], tmp31[117], tmp31[116], tmp31[115], tmp31[114], tmp31[113], tmp31[112], tmp31[111], tmp31[110], tmp31[109], tmp31[108], tmp31[107], tmp31[106], tmp31[105], tmp31[104], tmp31[103], tmp31[102], tmp31[101], tmp31[100], tmp31[99], tmp31[98], tmp31[97], tmp31[96], tmp31[95], tmp31[94], tmp31[93], tmp31[92], tmp31[91], tmp31[90], tmp31[89], tmp31[88], tmp31[87], tmp31[86], tmp31[85], tmp31[84], tmp31[83], tmp31[82], tmp31[81], tmp31[80], tmp31[79], tmp31[78], tmp31[77], tmp31[76], tmp31[75], tmp31[74], tmp31[73], tmp31[72], tmp31[71], tmp31[70], tmp31[69], tmp31[68], tmp31[67], tmp31[66], tmp31[65], tmp31[64], tmp31[63], tmp31[62], tmp31[61], tmp31[60], tmp31[59], tmp31[58], tmp31[57], tmp31[56], tmp31[55], tmp31[54], tmp31[53], tmp31[52], tmp31[51], tmp31[50], tmp31[49], tmp31[48], tmp31[47], tmp31[46], tmp31[45], tmp31[44], tmp31[43], tmp31[42], tmp31[41], tmp31[40], tmp31[39], tmp31[38], tmp31[37], tmp31[36], tmp31[35], tmp31[34], tmp31[33], tmp31[32], tmp31[31], tmp31[30], tmp31[29], tmp31[28], tmp31[27], tmp31[26], tmp31[25], tmp31[24], tmp31[23], tmp31[22], tmp31[21], tmp31[20], tmp31[19], tmp31[18], tmp31[17], tmp31[16], tmp31[15], tmp31[14], tmp31[13], tmp31[12], tmp31[11], tmp31[10], tmp31[9], tmp31[8], tmp31[7], tmp31[6], tmp31[5], tmp31[4], tmp31[3], tmp31[2], tmp31[1], tmp31[0]};
    assign tmp4997 = {tmp4996, const_447_0};
    assign tmp4998 = {const_448_0};
    assign tmp4999 = {tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998, tmp4998};
    assign tmp5000 = {tmp4999, const_448_0};
    assign tmp5001 = {tmp31[255]};
    assign tmp5002 = tmp5000 - tmp31;
    assign tmp5003 = {tmp5002[256]};
    assign tmp5004 = {tmp5000[255]};
    assign tmp5005 = ~tmp5004;
    assign tmp5006 = tmp5003 ^ tmp5005;
    assign tmp5007 = {tmp31[255]};
    assign tmp5008 = ~tmp5007;
    assign tmp5009 = tmp5006 ^ tmp5008;
    assign tmp5010 = {tmp4997[255]};
    assign tmp5011 = {const_449_0};
    assign tmp5012 = {tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011, tmp5011};
    assign tmp5013 = {tmp5012, const_449_0};
    assign tmp5014 = tmp4997 - tmp5013;
    assign tmp5015 = {tmp5014[256]};
    assign tmp5016 = {tmp4997[255]};
    assign tmp5017 = ~tmp5016;
    assign tmp5018 = tmp5015 ^ tmp5017;
    assign tmp5019 = {tmp5013[255]};
    assign tmp5020 = ~tmp5019;
    assign tmp5021 = tmp5018 ^ tmp5020;
    assign tmp5022 = tmp5009 & tmp5021;
    assign tmp5023 = {tmp31[255]};
    assign tmp5024 = {const_450_0};
    assign tmp5025 = {tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024, tmp5024};
    assign tmp5026 = {tmp5025, const_450_0};
    assign tmp5027 = tmp31 - tmp5026;
    assign tmp5028 = {tmp5027[256]};
    assign tmp5029 = {tmp31[255]};
    assign tmp5030 = ~tmp5029;
    assign tmp5031 = tmp5028 ^ tmp5030;
    assign tmp5032 = {tmp5026[255]};
    assign tmp5033 = ~tmp5032;
    assign tmp5034 = tmp5031 ^ tmp5033;
    assign tmp5035 = {const_451_0};
    assign tmp5036 = {tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035, tmp5035};
    assign tmp5037 = {tmp5036, const_451_0};
    assign tmp5038 = {tmp4997[255]};
    assign tmp5039 = tmp5037 - tmp4997;
    assign tmp5040 = {tmp5039[256]};
    assign tmp5041 = {tmp5037[255]};
    assign tmp5042 = ~tmp5041;
    assign tmp5043 = tmp5040 ^ tmp5042;
    assign tmp5044 = {tmp4997[255]};
    assign tmp5045 = ~tmp5044;
    assign tmp5046 = tmp5043 ^ tmp5045;
    assign tmp5047 = tmp5037 == tmp4997;
    assign tmp5048 = tmp5046 | tmp5047;
    assign tmp5049 = tmp5034 & tmp5048;
    assign tmp5050 = tmp5022 ? const_452_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp4997;
    assign tmp5051 = tmp5049 ? _ver_out_tmp_10 : tmp5050;
    assign tmp5052 = ~tmp35;
    assign tmp5053 = ~tmp36;
    assign tmp5054 = tmp5052 & tmp5053;
    assign tmp5055 = ~tmp57;
    assign tmp5056 = tmp5054 & tmp5055;
    assign tmp5057 = ~tmp1034;
    assign tmp5058 = tmp5056 & tmp5057;
    assign tmp5059 = tmp5058 & tmp2071;
    assign tmp5060 = ~tmp2583;
    assign tmp5061 = tmp5059 & tmp5060;
    assign tmp5062 = tmp5061 & tmp23;
    assign tmp5063 = ~tmp2627;
    assign tmp5064 = tmp5062 & tmp5063;
    assign tmp5065 = ~tmp2798;
    assign tmp5066 = tmp5064 & tmp5065;
    assign tmp5067 = ~tmp3425;
    assign tmp5068 = tmp5066 & tmp5067;
    assign tmp5069 = ~tmp4020;
    assign tmp5070 = tmp5068 & tmp5069;
    assign tmp5071 = tmp5070 & cfg_speculative_egest;
    assign tmp5072 = tmp5071 & tmp4511;
    assign tmp5073 = ~tmp24;
    assign tmp5074 = tmp5072 & tmp5073;
    assign tmp5075 = {tmp32[254], tmp32[253], tmp32[252], tmp32[251], tmp32[250], tmp32[249], tmp32[248], tmp32[247], tmp32[246], tmp32[245], tmp32[244], tmp32[243], tmp32[242], tmp32[241], tmp32[240], tmp32[239], tmp32[238], tmp32[237], tmp32[236], tmp32[235], tmp32[234], tmp32[233], tmp32[232], tmp32[231], tmp32[230], tmp32[229], tmp32[228], tmp32[227], tmp32[226], tmp32[225], tmp32[224], tmp32[223], tmp32[222], tmp32[221], tmp32[220], tmp32[219], tmp32[218], tmp32[217], tmp32[216], tmp32[215], tmp32[214], tmp32[213], tmp32[212], tmp32[211], tmp32[210], tmp32[209], tmp32[208], tmp32[207], tmp32[206], tmp32[205], tmp32[204], tmp32[203], tmp32[202], tmp32[201], tmp32[200], tmp32[199], tmp32[198], tmp32[197], tmp32[196], tmp32[195], tmp32[194], tmp32[193], tmp32[192], tmp32[191], tmp32[190], tmp32[189], tmp32[188], tmp32[187], tmp32[186], tmp32[185], tmp32[184], tmp32[183], tmp32[182], tmp32[181], tmp32[180], tmp32[179], tmp32[178], tmp32[177], tmp32[176], tmp32[175], tmp32[174], tmp32[173], tmp32[172], tmp32[171], tmp32[170], tmp32[169], tmp32[168], tmp32[167], tmp32[166], tmp32[165], tmp32[164], tmp32[163], tmp32[162], tmp32[161], tmp32[160], tmp32[159], tmp32[158], tmp32[157], tmp32[156], tmp32[155], tmp32[154], tmp32[153], tmp32[152], tmp32[151], tmp32[150], tmp32[149], tmp32[148], tmp32[147], tmp32[146], tmp32[145], tmp32[144], tmp32[143], tmp32[142], tmp32[141], tmp32[140], tmp32[139], tmp32[138], tmp32[137], tmp32[136], tmp32[135], tmp32[134], tmp32[133], tmp32[132], tmp32[131], tmp32[130], tmp32[129], tmp32[128], tmp32[127], tmp32[126], tmp32[125], tmp32[124], tmp32[123], tmp32[122], tmp32[121], tmp32[120], tmp32[119], tmp32[118], tmp32[117], tmp32[116], tmp32[115], tmp32[114], tmp32[113], tmp32[112], tmp32[111], tmp32[110], tmp32[109], tmp32[108], tmp32[107], tmp32[106], tmp32[105], tmp32[104], tmp32[103], tmp32[102], tmp32[101], tmp32[100], tmp32[99], tmp32[98], tmp32[97], tmp32[96], tmp32[95], tmp32[94], tmp32[93], tmp32[92], tmp32[91], tmp32[90], tmp32[89], tmp32[88], tmp32[87], tmp32[86], tmp32[85], tmp32[84], tmp32[83], tmp32[82], tmp32[81], tmp32[80], tmp32[79], tmp32[78], tmp32[77], tmp32[76], tmp32[75], tmp32[74], tmp32[73], tmp32[72], tmp32[71], tmp32[70], tmp32[69], tmp32[68], tmp32[67], tmp32[66], tmp32[65], tmp32[64], tmp32[63], tmp32[62], tmp32[61], tmp32[60], tmp32[59], tmp32[58], tmp32[57], tmp32[56], tmp32[55], tmp32[54], tmp32[53], tmp32[52], tmp32[51], tmp32[50], tmp32[49], tmp32[48], tmp32[47], tmp32[46], tmp32[45], tmp32[44], tmp32[43], tmp32[42], tmp32[41], tmp32[40], tmp32[39], tmp32[38], tmp32[37], tmp32[36], tmp32[35], tmp32[34], tmp32[33], tmp32[32], tmp32[31], tmp32[30], tmp32[29], tmp32[28], tmp32[27], tmp32[26], tmp32[25], tmp32[24], tmp32[23], tmp32[22], tmp32[21], tmp32[20], tmp32[19], tmp32[18], tmp32[17], tmp32[16], tmp32[15], tmp32[14], tmp32[13], tmp32[12], tmp32[11], tmp32[10], tmp32[9], tmp32[8], tmp32[7], tmp32[6], tmp32[5], tmp32[4], tmp32[3], tmp32[2], tmp32[1], tmp32[0]};
    assign tmp5076 = {tmp5075, const_454_0};
    assign tmp5077 = {const_455_0};
    assign tmp5078 = {tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077, tmp5077};
    assign tmp5079 = {tmp5078, const_455_0};
    assign tmp5080 = {tmp32[255]};
    assign tmp5081 = tmp5079 - tmp32;
    assign tmp5082 = {tmp5081[256]};
    assign tmp5083 = {tmp5079[255]};
    assign tmp5084 = ~tmp5083;
    assign tmp5085 = tmp5082 ^ tmp5084;
    assign tmp5086 = {tmp32[255]};
    assign tmp5087 = ~tmp5086;
    assign tmp5088 = tmp5085 ^ tmp5087;
    assign tmp5089 = {tmp5076[255]};
    assign tmp5090 = {const_456_0};
    assign tmp5091 = {tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090, tmp5090};
    assign tmp5092 = {tmp5091, const_456_0};
    assign tmp5093 = tmp5076 - tmp5092;
    assign tmp5094 = {tmp5093[256]};
    assign tmp5095 = {tmp5076[255]};
    assign tmp5096 = ~tmp5095;
    assign tmp5097 = tmp5094 ^ tmp5096;
    assign tmp5098 = {tmp5092[255]};
    assign tmp5099 = ~tmp5098;
    assign tmp5100 = tmp5097 ^ tmp5099;
    assign tmp5101 = tmp5088 & tmp5100;
    assign tmp5102 = {tmp32[255]};
    assign tmp5103 = {const_457_0};
    assign tmp5104 = {tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103, tmp5103};
    assign tmp5105 = {tmp5104, const_457_0};
    assign tmp5106 = tmp32 - tmp5105;
    assign tmp5107 = {tmp5106[256]};
    assign tmp5108 = {tmp32[255]};
    assign tmp5109 = ~tmp5108;
    assign tmp5110 = tmp5107 ^ tmp5109;
    assign tmp5111 = {tmp5105[255]};
    assign tmp5112 = ~tmp5111;
    assign tmp5113 = tmp5110 ^ tmp5112;
    assign tmp5114 = {const_458_0};
    assign tmp5115 = {tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114, tmp5114};
    assign tmp5116 = {tmp5115, const_458_0};
    assign tmp5117 = {tmp5076[255]};
    assign tmp5118 = tmp5116 - tmp5076;
    assign tmp5119 = {tmp5118[256]};
    assign tmp5120 = {tmp5116[255]};
    assign tmp5121 = ~tmp5120;
    assign tmp5122 = tmp5119 ^ tmp5121;
    assign tmp5123 = {tmp5076[255]};
    assign tmp5124 = ~tmp5123;
    assign tmp5125 = tmp5122 ^ tmp5124;
    assign tmp5126 = tmp5116 == tmp5076;
    assign tmp5127 = tmp5125 | tmp5126;
    assign tmp5128 = tmp5113 & tmp5127;
    assign tmp5129 = tmp5101 ? const_459_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp5076;
    assign tmp5130 = tmp5128 ? _ver_out_tmp_12 : tmp5129;
    assign tmp5131 = ~tmp35;
    assign tmp5132 = ~tmp36;
    assign tmp5133 = tmp5131 & tmp5132;
    assign tmp5134 = ~tmp57;
    assign tmp5135 = tmp5133 & tmp5134;
    assign tmp5136 = ~tmp1034;
    assign tmp5137 = tmp5135 & tmp5136;
    assign tmp5138 = tmp5137 & tmp2071;
    assign tmp5139 = ~tmp2583;
    assign tmp5140 = tmp5138 & tmp5139;
    assign tmp5141 = tmp5140 & tmp23;
    assign tmp5142 = ~tmp2627;
    assign tmp5143 = tmp5141 & tmp5142;
    assign tmp5144 = ~tmp2798;
    assign tmp5145 = tmp5143 & tmp5144;
    assign tmp5146 = ~tmp3425;
    assign tmp5147 = tmp5145 & tmp5146;
    assign tmp5148 = ~tmp4020;
    assign tmp5149 = tmp5147 & tmp5148;
    assign tmp5150 = tmp5149 & cfg_speculative_egest;
    assign tmp5151 = tmp5150 & tmp4511;
    assign tmp5152 = ~tmp24;
    assign tmp5153 = tmp5151 & tmp5152;
    assign tmp5154 = {tmp25[254], tmp25[253], tmp25[252], tmp25[251], tmp25[250], tmp25[249], tmp25[248], tmp25[247], tmp25[246], tmp25[245], tmp25[244], tmp25[243], tmp25[242], tmp25[241], tmp25[240], tmp25[239], tmp25[238], tmp25[237], tmp25[236], tmp25[235], tmp25[234], tmp25[233], tmp25[232], tmp25[231], tmp25[230], tmp25[229], tmp25[228], tmp25[227], tmp25[226], tmp25[225], tmp25[224], tmp25[223], tmp25[222], tmp25[221], tmp25[220], tmp25[219], tmp25[218], tmp25[217], tmp25[216], tmp25[215], tmp25[214], tmp25[213], tmp25[212], tmp25[211], tmp25[210], tmp25[209], tmp25[208], tmp25[207], tmp25[206], tmp25[205], tmp25[204], tmp25[203], tmp25[202], tmp25[201], tmp25[200], tmp25[199], tmp25[198], tmp25[197], tmp25[196], tmp25[195], tmp25[194], tmp25[193], tmp25[192], tmp25[191], tmp25[190], tmp25[189], tmp25[188], tmp25[187], tmp25[186], tmp25[185], tmp25[184], tmp25[183], tmp25[182], tmp25[181], tmp25[180], tmp25[179], tmp25[178], tmp25[177], tmp25[176], tmp25[175], tmp25[174], tmp25[173], tmp25[172], tmp25[171], tmp25[170], tmp25[169], tmp25[168], tmp25[167], tmp25[166], tmp25[165], tmp25[164], tmp25[163], tmp25[162], tmp25[161], tmp25[160], tmp25[159], tmp25[158], tmp25[157], tmp25[156], tmp25[155], tmp25[154], tmp25[153], tmp25[152], tmp25[151], tmp25[150], tmp25[149], tmp25[148], tmp25[147], tmp25[146], tmp25[145], tmp25[144], tmp25[143], tmp25[142], tmp25[141], tmp25[140], tmp25[139], tmp25[138], tmp25[137], tmp25[136], tmp25[135], tmp25[134], tmp25[133], tmp25[132], tmp25[131], tmp25[130], tmp25[129], tmp25[128], tmp25[127], tmp25[126], tmp25[125], tmp25[124], tmp25[123], tmp25[122], tmp25[121], tmp25[120], tmp25[119], tmp25[118], tmp25[117], tmp25[116], tmp25[115], tmp25[114], tmp25[113], tmp25[112], tmp25[111], tmp25[110], tmp25[109], tmp25[108], tmp25[107], tmp25[106], tmp25[105], tmp25[104], tmp25[103], tmp25[102], tmp25[101], tmp25[100], tmp25[99], tmp25[98], tmp25[97], tmp25[96], tmp25[95], tmp25[94], tmp25[93], tmp25[92], tmp25[91], tmp25[90], tmp25[89], tmp25[88], tmp25[87], tmp25[86], tmp25[85], tmp25[84], tmp25[83], tmp25[82], tmp25[81], tmp25[80], tmp25[79], tmp25[78], tmp25[77], tmp25[76], tmp25[75], tmp25[74], tmp25[73], tmp25[72], tmp25[71], tmp25[70], tmp25[69], tmp25[68], tmp25[67], tmp25[66], tmp25[65], tmp25[64], tmp25[63], tmp25[62], tmp25[61], tmp25[60], tmp25[59], tmp25[58], tmp25[57], tmp25[56], tmp25[55], tmp25[54], tmp25[53], tmp25[52], tmp25[51], tmp25[50], tmp25[49], tmp25[48], tmp25[47], tmp25[46], tmp25[45], tmp25[44], tmp25[43], tmp25[42], tmp25[41], tmp25[40], tmp25[39], tmp25[38], tmp25[37], tmp25[36], tmp25[35], tmp25[34], tmp25[33], tmp25[32], tmp25[31], tmp25[30], tmp25[29], tmp25[28], tmp25[27], tmp25[26], tmp25[25], tmp25[24], tmp25[23], tmp25[22], tmp25[21], tmp25[20], tmp25[19], tmp25[18], tmp25[17], tmp25[16], tmp25[15], tmp25[14], tmp25[13], tmp25[12], tmp25[11], tmp25[10], tmp25[9], tmp25[8], tmp25[7], tmp25[6], tmp25[5], tmp25[4], tmp25[3], tmp25[2], tmp25[1], tmp25[0]};
    assign tmp5155 = {tmp5154, const_461_0};
    assign tmp5156 = {const_462_0};
    assign tmp5157 = {tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156, tmp5156};
    assign tmp5158 = {tmp5157, const_462_0};
    assign tmp5159 = {tmp25[255]};
    assign tmp5160 = tmp5158 - tmp25;
    assign tmp5161 = {tmp5160[256]};
    assign tmp5162 = {tmp5158[255]};
    assign tmp5163 = ~tmp5162;
    assign tmp5164 = tmp5161 ^ tmp5163;
    assign tmp5165 = {tmp25[255]};
    assign tmp5166 = ~tmp5165;
    assign tmp5167 = tmp5164 ^ tmp5166;
    assign tmp5168 = {tmp5155[255]};
    assign tmp5169 = {const_463_0};
    assign tmp5170 = {tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169, tmp5169};
    assign tmp5171 = {tmp5170, const_463_0};
    assign tmp5172 = tmp5155 - tmp5171;
    assign tmp5173 = {tmp5172[256]};
    assign tmp5174 = {tmp5155[255]};
    assign tmp5175 = ~tmp5174;
    assign tmp5176 = tmp5173 ^ tmp5175;
    assign tmp5177 = {tmp5171[255]};
    assign tmp5178 = ~tmp5177;
    assign tmp5179 = tmp5176 ^ tmp5178;
    assign tmp5180 = tmp5167 & tmp5179;
    assign tmp5181 = {tmp25[255]};
    assign tmp5182 = {const_464_0};
    assign tmp5183 = {tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182, tmp5182};
    assign tmp5184 = {tmp5183, const_464_0};
    assign tmp5185 = tmp25 - tmp5184;
    assign tmp5186 = {tmp5185[256]};
    assign tmp5187 = {tmp25[255]};
    assign tmp5188 = ~tmp5187;
    assign tmp5189 = tmp5186 ^ tmp5188;
    assign tmp5190 = {tmp5184[255]};
    assign tmp5191 = ~tmp5190;
    assign tmp5192 = tmp5189 ^ tmp5191;
    assign tmp5193 = {const_465_0};
    assign tmp5194 = {tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193, tmp5193};
    assign tmp5195 = {tmp5194, const_465_0};
    assign tmp5196 = {tmp5155[255]};
    assign tmp5197 = tmp5195 - tmp5155;
    assign tmp5198 = {tmp5197[256]};
    assign tmp5199 = {tmp5195[255]};
    assign tmp5200 = ~tmp5199;
    assign tmp5201 = tmp5198 ^ tmp5200;
    assign tmp5202 = {tmp5155[255]};
    assign tmp5203 = ~tmp5202;
    assign tmp5204 = tmp5201 ^ tmp5203;
    assign tmp5205 = tmp5195 == tmp5155;
    assign tmp5206 = tmp5204 | tmp5205;
    assign tmp5207 = tmp5192 & tmp5206;
    assign tmp5208 = tmp5180 ? const_466_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp5155;
    assign tmp5209 = tmp5207 ? _ver_out_tmp_14 : tmp5208;
    assign tmp5210 = {tmp29[255]};
    assign tmp5211 = {tmp5209[255]};
    assign tmp5212 = tmp29 - tmp5209;
    assign tmp5213 = {tmp5212[256]};
    assign tmp5214 = {tmp29[255]};
    assign tmp5215 = ~tmp5214;
    assign tmp5216 = tmp5213 ^ tmp5215;
    assign tmp5217 = {tmp5209[255]};
    assign tmp5218 = ~tmp5217;
    assign tmp5219 = tmp5216 ^ tmp5218;
    assign tmp5220 = {tmp29[254], tmp29[253], tmp29[252], tmp29[251], tmp29[250], tmp29[249], tmp29[248], tmp29[247], tmp29[246], tmp29[245], tmp29[244], tmp29[243], tmp29[242], tmp29[241], tmp29[240], tmp29[239], tmp29[238], tmp29[237], tmp29[236], tmp29[235], tmp29[234], tmp29[233], tmp29[232], tmp29[231], tmp29[230], tmp29[229], tmp29[228], tmp29[227], tmp29[226], tmp29[225], tmp29[224], tmp29[223], tmp29[222], tmp29[221], tmp29[220], tmp29[219], tmp29[218], tmp29[217], tmp29[216], tmp29[215], tmp29[214], tmp29[213], tmp29[212], tmp29[211], tmp29[210], tmp29[209], tmp29[208], tmp29[207], tmp29[206], tmp29[205], tmp29[204], tmp29[203], tmp29[202], tmp29[201], tmp29[200], tmp29[199], tmp29[198], tmp29[197], tmp29[196], tmp29[195], tmp29[194], tmp29[193], tmp29[192], tmp29[191], tmp29[190], tmp29[189], tmp29[188], tmp29[187], tmp29[186], tmp29[185], tmp29[184], tmp29[183], tmp29[182], tmp29[181], tmp29[180], tmp29[179], tmp29[178], tmp29[177], tmp29[176], tmp29[175], tmp29[174], tmp29[173], tmp29[172], tmp29[171], tmp29[170], tmp29[169], tmp29[168], tmp29[167], tmp29[166], tmp29[165], tmp29[164], tmp29[163], tmp29[162], tmp29[161], tmp29[160], tmp29[159], tmp29[158], tmp29[157], tmp29[156], tmp29[155], tmp29[154], tmp29[153], tmp29[152], tmp29[151], tmp29[150], tmp29[149], tmp29[148], tmp29[147], tmp29[146], tmp29[145], tmp29[144], tmp29[143], tmp29[142], tmp29[141], tmp29[140], tmp29[139], tmp29[138], tmp29[137], tmp29[136], tmp29[135], tmp29[134], tmp29[133], tmp29[132], tmp29[131], tmp29[130], tmp29[129], tmp29[128], tmp29[127], tmp29[126], tmp29[125], tmp29[124], tmp29[123], tmp29[122], tmp29[121], tmp29[120], tmp29[119], tmp29[118], tmp29[117], tmp29[116], tmp29[115], tmp29[114], tmp29[113], tmp29[112], tmp29[111], tmp29[110], tmp29[109], tmp29[108], tmp29[107], tmp29[106], tmp29[105], tmp29[104], tmp29[103], tmp29[102], tmp29[101], tmp29[100], tmp29[99], tmp29[98], tmp29[97], tmp29[96], tmp29[95], tmp29[94], tmp29[93], tmp29[92], tmp29[91], tmp29[90], tmp29[89], tmp29[88], tmp29[87], tmp29[86], tmp29[85], tmp29[84], tmp29[83], tmp29[82], tmp29[81], tmp29[80], tmp29[79], tmp29[78], tmp29[77], tmp29[76], tmp29[75], tmp29[74], tmp29[73], tmp29[72], tmp29[71], tmp29[70], tmp29[69], tmp29[68], tmp29[67], tmp29[66], tmp29[65], tmp29[64], tmp29[63], tmp29[62], tmp29[61], tmp29[60], tmp29[59], tmp29[58], tmp29[57], tmp29[56], tmp29[55], tmp29[54], tmp29[53], tmp29[52], tmp29[51], tmp29[50], tmp29[49], tmp29[48], tmp29[47], tmp29[46], tmp29[45], tmp29[44], tmp29[43], tmp29[42], tmp29[41], tmp29[40], tmp29[39], tmp29[38], tmp29[37], tmp29[36], tmp29[35], tmp29[34], tmp29[33], tmp29[32], tmp29[31], tmp29[30], tmp29[29], tmp29[28], tmp29[27], tmp29[26], tmp29[25], tmp29[24], tmp29[23], tmp29[22], tmp29[21], tmp29[20], tmp29[19], tmp29[18], tmp29[17], tmp29[16], tmp29[15], tmp29[14], tmp29[13], tmp29[12], tmp29[11], tmp29[10], tmp29[9], tmp29[8], tmp29[7], tmp29[6], tmp29[5], tmp29[4], tmp29[3], tmp29[2], tmp29[1], tmp29[0]};
    assign tmp5221 = {tmp5220, const_468_0};
    assign tmp5222 = {const_469_0};
    assign tmp5223 = {tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222, tmp5222};
    assign tmp5224 = {tmp5223, const_469_0};
    assign tmp5225 = {tmp29[255]};
    assign tmp5226 = tmp5224 - tmp29;
    assign tmp5227 = {tmp5226[256]};
    assign tmp5228 = {tmp5224[255]};
    assign tmp5229 = ~tmp5228;
    assign tmp5230 = tmp5227 ^ tmp5229;
    assign tmp5231 = {tmp29[255]};
    assign tmp5232 = ~tmp5231;
    assign tmp5233 = tmp5230 ^ tmp5232;
    assign tmp5234 = {tmp5221[255]};
    assign tmp5235 = {const_470_0};
    assign tmp5236 = {tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235, tmp5235};
    assign tmp5237 = {tmp5236, const_470_0};
    assign tmp5238 = tmp5221 - tmp5237;
    assign tmp5239 = {tmp5238[256]};
    assign tmp5240 = {tmp5221[255]};
    assign tmp5241 = ~tmp5240;
    assign tmp5242 = tmp5239 ^ tmp5241;
    assign tmp5243 = {tmp5237[255]};
    assign tmp5244 = ~tmp5243;
    assign tmp5245 = tmp5242 ^ tmp5244;
    assign tmp5246 = tmp5233 & tmp5245;
    assign tmp5247 = {tmp29[255]};
    assign tmp5248 = {const_471_0};
    assign tmp5249 = {tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248, tmp5248};
    assign tmp5250 = {tmp5249, const_471_0};
    assign tmp5251 = tmp29 - tmp5250;
    assign tmp5252 = {tmp5251[256]};
    assign tmp5253 = {tmp29[255]};
    assign tmp5254 = ~tmp5253;
    assign tmp5255 = tmp5252 ^ tmp5254;
    assign tmp5256 = {tmp5250[255]};
    assign tmp5257 = ~tmp5256;
    assign tmp5258 = tmp5255 ^ tmp5257;
    assign tmp5259 = {const_472_0};
    assign tmp5260 = {tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259, tmp5259};
    assign tmp5261 = {tmp5260, const_472_0};
    assign tmp5262 = {tmp5221[255]};
    assign tmp5263 = tmp5261 - tmp5221;
    assign tmp5264 = {tmp5263[256]};
    assign tmp5265 = {tmp5261[255]};
    assign tmp5266 = ~tmp5265;
    assign tmp5267 = tmp5264 ^ tmp5266;
    assign tmp5268 = {tmp5221[255]};
    assign tmp5269 = ~tmp5268;
    assign tmp5270 = tmp5267 ^ tmp5269;
    assign tmp5271 = tmp5261 == tmp5221;
    assign tmp5272 = tmp5270 | tmp5271;
    assign tmp5273 = tmp5258 & tmp5272;
    assign tmp5274 = tmp5246 ? const_473_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp5221;
    assign tmp5275 = tmp5273 ? _ver_out_tmp_18 : tmp5274;
    assign tmp5276 = {tmp25[255]};
    assign tmp5277 = {tmp5275[255]};
    assign tmp5278 = tmp25 - tmp5275;
    assign tmp5279 = {tmp5278[256]};
    assign tmp5280 = {tmp25[255]};
    assign tmp5281 = ~tmp5280;
    assign tmp5282 = tmp5279 ^ tmp5281;
    assign tmp5283 = {tmp5275[255]};
    assign tmp5284 = ~tmp5283;
    assign tmp5285 = tmp5282 ^ tmp5284;
    assign tmp5286 = tmp5219 & tmp5285;
    assign tmp5287 = {tmp26[254], tmp26[253], tmp26[252], tmp26[251], tmp26[250], tmp26[249], tmp26[248], tmp26[247], tmp26[246], tmp26[245], tmp26[244], tmp26[243], tmp26[242], tmp26[241], tmp26[240], tmp26[239], tmp26[238], tmp26[237], tmp26[236], tmp26[235], tmp26[234], tmp26[233], tmp26[232], tmp26[231], tmp26[230], tmp26[229], tmp26[228], tmp26[227], tmp26[226], tmp26[225], tmp26[224], tmp26[223], tmp26[222], tmp26[221], tmp26[220], tmp26[219], tmp26[218], tmp26[217], tmp26[216], tmp26[215], tmp26[214], tmp26[213], tmp26[212], tmp26[211], tmp26[210], tmp26[209], tmp26[208], tmp26[207], tmp26[206], tmp26[205], tmp26[204], tmp26[203], tmp26[202], tmp26[201], tmp26[200], tmp26[199], tmp26[198], tmp26[197], tmp26[196], tmp26[195], tmp26[194], tmp26[193], tmp26[192], tmp26[191], tmp26[190], tmp26[189], tmp26[188], tmp26[187], tmp26[186], tmp26[185], tmp26[184], tmp26[183], tmp26[182], tmp26[181], tmp26[180], tmp26[179], tmp26[178], tmp26[177], tmp26[176], tmp26[175], tmp26[174], tmp26[173], tmp26[172], tmp26[171], tmp26[170], tmp26[169], tmp26[168], tmp26[167], tmp26[166], tmp26[165], tmp26[164], tmp26[163], tmp26[162], tmp26[161], tmp26[160], tmp26[159], tmp26[158], tmp26[157], tmp26[156], tmp26[155], tmp26[154], tmp26[153], tmp26[152], tmp26[151], tmp26[150], tmp26[149], tmp26[148], tmp26[147], tmp26[146], tmp26[145], tmp26[144], tmp26[143], tmp26[142], tmp26[141], tmp26[140], tmp26[139], tmp26[138], tmp26[137], tmp26[136], tmp26[135], tmp26[134], tmp26[133], tmp26[132], tmp26[131], tmp26[130], tmp26[129], tmp26[128], tmp26[127], tmp26[126], tmp26[125], tmp26[124], tmp26[123], tmp26[122], tmp26[121], tmp26[120], tmp26[119], tmp26[118], tmp26[117], tmp26[116], tmp26[115], tmp26[114], tmp26[113], tmp26[112], tmp26[111], tmp26[110], tmp26[109], tmp26[108], tmp26[107], tmp26[106], tmp26[105], tmp26[104], tmp26[103], tmp26[102], tmp26[101], tmp26[100], tmp26[99], tmp26[98], tmp26[97], tmp26[96], tmp26[95], tmp26[94], tmp26[93], tmp26[92], tmp26[91], tmp26[90], tmp26[89], tmp26[88], tmp26[87], tmp26[86], tmp26[85], tmp26[84], tmp26[83], tmp26[82], tmp26[81], tmp26[80], tmp26[79], tmp26[78], tmp26[77], tmp26[76], tmp26[75], tmp26[74], tmp26[73], tmp26[72], tmp26[71], tmp26[70], tmp26[69], tmp26[68], tmp26[67], tmp26[66], tmp26[65], tmp26[64], tmp26[63], tmp26[62], tmp26[61], tmp26[60], tmp26[59], tmp26[58], tmp26[57], tmp26[56], tmp26[55], tmp26[54], tmp26[53], tmp26[52], tmp26[51], tmp26[50], tmp26[49], tmp26[48], tmp26[47], tmp26[46], tmp26[45], tmp26[44], tmp26[43], tmp26[42], tmp26[41], tmp26[40], tmp26[39], tmp26[38], tmp26[37], tmp26[36], tmp26[35], tmp26[34], tmp26[33], tmp26[32], tmp26[31], tmp26[30], tmp26[29], tmp26[28], tmp26[27], tmp26[26], tmp26[25], tmp26[24], tmp26[23], tmp26[22], tmp26[21], tmp26[20], tmp26[19], tmp26[18], tmp26[17], tmp26[16], tmp26[15], tmp26[14], tmp26[13], tmp26[12], tmp26[11], tmp26[10], tmp26[9], tmp26[8], tmp26[7], tmp26[6], tmp26[5], tmp26[4], tmp26[3], tmp26[2], tmp26[1], tmp26[0]};
    assign tmp5288 = {tmp5287, const_475_0};
    assign tmp5289 = {const_476_0};
    assign tmp5290 = {tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289, tmp5289};
    assign tmp5291 = {tmp5290, const_476_0};
    assign tmp5292 = {tmp26[255]};
    assign tmp5293 = tmp5291 - tmp26;
    assign tmp5294 = {tmp5293[256]};
    assign tmp5295 = {tmp5291[255]};
    assign tmp5296 = ~tmp5295;
    assign tmp5297 = tmp5294 ^ tmp5296;
    assign tmp5298 = {tmp26[255]};
    assign tmp5299 = ~tmp5298;
    assign tmp5300 = tmp5297 ^ tmp5299;
    assign tmp5301 = {tmp5288[255]};
    assign tmp5302 = {const_477_0};
    assign tmp5303 = {tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302, tmp5302};
    assign tmp5304 = {tmp5303, const_477_0};
    assign tmp5305 = tmp5288 - tmp5304;
    assign tmp5306 = {tmp5305[256]};
    assign tmp5307 = {tmp5288[255]};
    assign tmp5308 = ~tmp5307;
    assign tmp5309 = tmp5306 ^ tmp5308;
    assign tmp5310 = {tmp5304[255]};
    assign tmp5311 = ~tmp5310;
    assign tmp5312 = tmp5309 ^ tmp5311;
    assign tmp5313 = tmp5300 & tmp5312;
    assign tmp5314 = {tmp26[255]};
    assign tmp5315 = {const_478_0};
    assign tmp5316 = {tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315, tmp5315};
    assign tmp5317 = {tmp5316, const_478_0};
    assign tmp5318 = tmp26 - tmp5317;
    assign tmp5319 = {tmp5318[256]};
    assign tmp5320 = {tmp26[255]};
    assign tmp5321 = ~tmp5320;
    assign tmp5322 = tmp5319 ^ tmp5321;
    assign tmp5323 = {tmp5317[255]};
    assign tmp5324 = ~tmp5323;
    assign tmp5325 = tmp5322 ^ tmp5324;
    assign tmp5326 = {const_479_0};
    assign tmp5327 = {tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326, tmp5326};
    assign tmp5328 = {tmp5327, const_479_0};
    assign tmp5329 = {tmp5288[255]};
    assign tmp5330 = tmp5328 - tmp5288;
    assign tmp5331 = {tmp5330[256]};
    assign tmp5332 = {tmp5328[255]};
    assign tmp5333 = ~tmp5332;
    assign tmp5334 = tmp5331 ^ tmp5333;
    assign tmp5335 = {tmp5288[255]};
    assign tmp5336 = ~tmp5335;
    assign tmp5337 = tmp5334 ^ tmp5336;
    assign tmp5338 = tmp5328 == tmp5288;
    assign tmp5339 = tmp5337 | tmp5338;
    assign tmp5340 = tmp5325 & tmp5339;
    assign tmp5341 = tmp5313 ? const_480_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp5288;
    assign tmp5342 = tmp5340 ? _ver_out_tmp_21 : tmp5341;
    assign tmp5343 = {tmp30[255]};
    assign tmp5344 = {tmp5342[255]};
    assign tmp5345 = tmp30 - tmp5342;
    assign tmp5346 = {tmp5345[256]};
    assign tmp5347 = {tmp30[255]};
    assign tmp5348 = ~tmp5347;
    assign tmp5349 = tmp5346 ^ tmp5348;
    assign tmp5350 = {tmp5342[255]};
    assign tmp5351 = ~tmp5350;
    assign tmp5352 = tmp5349 ^ tmp5351;
    assign tmp5353 = tmp5286 & tmp5352;
    assign tmp5354 = {tmp30[254], tmp30[253], tmp30[252], tmp30[251], tmp30[250], tmp30[249], tmp30[248], tmp30[247], tmp30[246], tmp30[245], tmp30[244], tmp30[243], tmp30[242], tmp30[241], tmp30[240], tmp30[239], tmp30[238], tmp30[237], tmp30[236], tmp30[235], tmp30[234], tmp30[233], tmp30[232], tmp30[231], tmp30[230], tmp30[229], tmp30[228], tmp30[227], tmp30[226], tmp30[225], tmp30[224], tmp30[223], tmp30[222], tmp30[221], tmp30[220], tmp30[219], tmp30[218], tmp30[217], tmp30[216], tmp30[215], tmp30[214], tmp30[213], tmp30[212], tmp30[211], tmp30[210], tmp30[209], tmp30[208], tmp30[207], tmp30[206], tmp30[205], tmp30[204], tmp30[203], tmp30[202], tmp30[201], tmp30[200], tmp30[199], tmp30[198], tmp30[197], tmp30[196], tmp30[195], tmp30[194], tmp30[193], tmp30[192], tmp30[191], tmp30[190], tmp30[189], tmp30[188], tmp30[187], tmp30[186], tmp30[185], tmp30[184], tmp30[183], tmp30[182], tmp30[181], tmp30[180], tmp30[179], tmp30[178], tmp30[177], tmp30[176], tmp30[175], tmp30[174], tmp30[173], tmp30[172], tmp30[171], tmp30[170], tmp30[169], tmp30[168], tmp30[167], tmp30[166], tmp30[165], tmp30[164], tmp30[163], tmp30[162], tmp30[161], tmp30[160], tmp30[159], tmp30[158], tmp30[157], tmp30[156], tmp30[155], tmp30[154], tmp30[153], tmp30[152], tmp30[151], tmp30[150], tmp30[149], tmp30[148], tmp30[147], tmp30[146], tmp30[145], tmp30[144], tmp30[143], tmp30[142], tmp30[141], tmp30[140], tmp30[139], tmp30[138], tmp30[137], tmp30[136], tmp30[135], tmp30[134], tmp30[133], tmp30[132], tmp30[131], tmp30[130], tmp30[129], tmp30[128], tmp30[127], tmp30[126], tmp30[125], tmp30[124], tmp30[123], tmp30[122], tmp30[121], tmp30[120], tmp30[119], tmp30[118], tmp30[117], tmp30[116], tmp30[115], tmp30[114], tmp30[113], tmp30[112], tmp30[111], tmp30[110], tmp30[109], tmp30[108], tmp30[107], tmp30[106], tmp30[105], tmp30[104], tmp30[103], tmp30[102], tmp30[101], tmp30[100], tmp30[99], tmp30[98], tmp30[97], tmp30[96], tmp30[95], tmp30[94], tmp30[93], tmp30[92], tmp30[91], tmp30[90], tmp30[89], tmp30[88], tmp30[87], tmp30[86], tmp30[85], tmp30[84], tmp30[83], tmp30[82], tmp30[81], tmp30[80], tmp30[79], tmp30[78], tmp30[77], tmp30[76], tmp30[75], tmp30[74], tmp30[73], tmp30[72], tmp30[71], tmp30[70], tmp30[69], tmp30[68], tmp30[67], tmp30[66], tmp30[65], tmp30[64], tmp30[63], tmp30[62], tmp30[61], tmp30[60], tmp30[59], tmp30[58], tmp30[57], tmp30[56], tmp30[55], tmp30[54], tmp30[53], tmp30[52], tmp30[51], tmp30[50], tmp30[49], tmp30[48], tmp30[47], tmp30[46], tmp30[45], tmp30[44], tmp30[43], tmp30[42], tmp30[41], tmp30[40], tmp30[39], tmp30[38], tmp30[37], tmp30[36], tmp30[35], tmp30[34], tmp30[33], tmp30[32], tmp30[31], tmp30[30], tmp30[29], tmp30[28], tmp30[27], tmp30[26], tmp30[25], tmp30[24], tmp30[23], tmp30[22], tmp30[21], tmp30[20], tmp30[19], tmp30[18], tmp30[17], tmp30[16], tmp30[15], tmp30[14], tmp30[13], tmp30[12], tmp30[11], tmp30[10], tmp30[9], tmp30[8], tmp30[7], tmp30[6], tmp30[5], tmp30[4], tmp30[3], tmp30[2], tmp30[1], tmp30[0]};
    assign tmp5355 = {tmp5354, const_482_0};
    assign tmp5356 = {const_483_0};
    assign tmp5357 = {tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356, tmp5356};
    assign tmp5358 = {tmp5357, const_483_0};
    assign tmp5359 = {tmp30[255]};
    assign tmp5360 = tmp5358 - tmp30;
    assign tmp5361 = {tmp5360[256]};
    assign tmp5362 = {tmp5358[255]};
    assign tmp5363 = ~tmp5362;
    assign tmp5364 = tmp5361 ^ tmp5363;
    assign tmp5365 = {tmp30[255]};
    assign tmp5366 = ~tmp5365;
    assign tmp5367 = tmp5364 ^ tmp5366;
    assign tmp5368 = {tmp5355[255]};
    assign tmp5369 = {const_484_0};
    assign tmp5370 = {tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369, tmp5369};
    assign tmp5371 = {tmp5370, const_484_0};
    assign tmp5372 = tmp5355 - tmp5371;
    assign tmp5373 = {tmp5372[256]};
    assign tmp5374 = {tmp5355[255]};
    assign tmp5375 = ~tmp5374;
    assign tmp5376 = tmp5373 ^ tmp5375;
    assign tmp5377 = {tmp5371[255]};
    assign tmp5378 = ~tmp5377;
    assign tmp5379 = tmp5376 ^ tmp5378;
    assign tmp5380 = tmp5367 & tmp5379;
    assign tmp5381 = {tmp30[255]};
    assign tmp5382 = {const_485_0};
    assign tmp5383 = {tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382, tmp5382};
    assign tmp5384 = {tmp5383, const_485_0};
    assign tmp5385 = tmp30 - tmp5384;
    assign tmp5386 = {tmp5385[256]};
    assign tmp5387 = {tmp30[255]};
    assign tmp5388 = ~tmp5387;
    assign tmp5389 = tmp5386 ^ tmp5388;
    assign tmp5390 = {tmp5384[255]};
    assign tmp5391 = ~tmp5390;
    assign tmp5392 = tmp5389 ^ tmp5391;
    assign tmp5393 = {const_486_0};
    assign tmp5394 = {tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393, tmp5393};
    assign tmp5395 = {tmp5394, const_486_0};
    assign tmp5396 = {tmp5355[255]};
    assign tmp5397 = tmp5395 - tmp5355;
    assign tmp5398 = {tmp5397[256]};
    assign tmp5399 = {tmp5395[255]};
    assign tmp5400 = ~tmp5399;
    assign tmp5401 = tmp5398 ^ tmp5400;
    assign tmp5402 = {tmp5355[255]};
    assign tmp5403 = ~tmp5402;
    assign tmp5404 = tmp5401 ^ tmp5403;
    assign tmp5405 = tmp5395 == tmp5355;
    assign tmp5406 = tmp5404 | tmp5405;
    assign tmp5407 = tmp5392 & tmp5406;
    assign tmp5408 = tmp5380 ? const_487_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp5355;
    assign tmp5409 = tmp5407 ? _ver_out_tmp_34 : tmp5408;
    assign tmp5410 = {tmp26[255]};
    assign tmp5411 = {tmp5409[255]};
    assign tmp5412 = tmp26 - tmp5409;
    assign tmp5413 = {tmp5412[256]};
    assign tmp5414 = {tmp26[255]};
    assign tmp5415 = ~tmp5414;
    assign tmp5416 = tmp5413 ^ tmp5415;
    assign tmp5417 = {tmp5409[255]};
    assign tmp5418 = ~tmp5417;
    assign tmp5419 = tmp5416 ^ tmp5418;
    assign tmp5420 = tmp5353 & tmp5419;
    assign tmp5421 = {tmp27[254], tmp27[253], tmp27[252], tmp27[251], tmp27[250], tmp27[249], tmp27[248], tmp27[247], tmp27[246], tmp27[245], tmp27[244], tmp27[243], tmp27[242], tmp27[241], tmp27[240], tmp27[239], tmp27[238], tmp27[237], tmp27[236], tmp27[235], tmp27[234], tmp27[233], tmp27[232], tmp27[231], tmp27[230], tmp27[229], tmp27[228], tmp27[227], tmp27[226], tmp27[225], tmp27[224], tmp27[223], tmp27[222], tmp27[221], tmp27[220], tmp27[219], tmp27[218], tmp27[217], tmp27[216], tmp27[215], tmp27[214], tmp27[213], tmp27[212], tmp27[211], tmp27[210], tmp27[209], tmp27[208], tmp27[207], tmp27[206], tmp27[205], tmp27[204], tmp27[203], tmp27[202], tmp27[201], tmp27[200], tmp27[199], tmp27[198], tmp27[197], tmp27[196], tmp27[195], tmp27[194], tmp27[193], tmp27[192], tmp27[191], tmp27[190], tmp27[189], tmp27[188], tmp27[187], tmp27[186], tmp27[185], tmp27[184], tmp27[183], tmp27[182], tmp27[181], tmp27[180], tmp27[179], tmp27[178], tmp27[177], tmp27[176], tmp27[175], tmp27[174], tmp27[173], tmp27[172], tmp27[171], tmp27[170], tmp27[169], tmp27[168], tmp27[167], tmp27[166], tmp27[165], tmp27[164], tmp27[163], tmp27[162], tmp27[161], tmp27[160], tmp27[159], tmp27[158], tmp27[157], tmp27[156], tmp27[155], tmp27[154], tmp27[153], tmp27[152], tmp27[151], tmp27[150], tmp27[149], tmp27[148], tmp27[147], tmp27[146], tmp27[145], tmp27[144], tmp27[143], tmp27[142], tmp27[141], tmp27[140], tmp27[139], tmp27[138], tmp27[137], tmp27[136], tmp27[135], tmp27[134], tmp27[133], tmp27[132], tmp27[131], tmp27[130], tmp27[129], tmp27[128], tmp27[127], tmp27[126], tmp27[125], tmp27[124], tmp27[123], tmp27[122], tmp27[121], tmp27[120], tmp27[119], tmp27[118], tmp27[117], tmp27[116], tmp27[115], tmp27[114], tmp27[113], tmp27[112], tmp27[111], tmp27[110], tmp27[109], tmp27[108], tmp27[107], tmp27[106], tmp27[105], tmp27[104], tmp27[103], tmp27[102], tmp27[101], tmp27[100], tmp27[99], tmp27[98], tmp27[97], tmp27[96], tmp27[95], tmp27[94], tmp27[93], tmp27[92], tmp27[91], tmp27[90], tmp27[89], tmp27[88], tmp27[87], tmp27[86], tmp27[85], tmp27[84], tmp27[83], tmp27[82], tmp27[81], tmp27[80], tmp27[79], tmp27[78], tmp27[77], tmp27[76], tmp27[75], tmp27[74], tmp27[73], tmp27[72], tmp27[71], tmp27[70], tmp27[69], tmp27[68], tmp27[67], tmp27[66], tmp27[65], tmp27[64], tmp27[63], tmp27[62], tmp27[61], tmp27[60], tmp27[59], tmp27[58], tmp27[57], tmp27[56], tmp27[55], tmp27[54], tmp27[53], tmp27[52], tmp27[51], tmp27[50], tmp27[49], tmp27[48], tmp27[47], tmp27[46], tmp27[45], tmp27[44], tmp27[43], tmp27[42], tmp27[41], tmp27[40], tmp27[39], tmp27[38], tmp27[37], tmp27[36], tmp27[35], tmp27[34], tmp27[33], tmp27[32], tmp27[31], tmp27[30], tmp27[29], tmp27[28], tmp27[27], tmp27[26], tmp27[25], tmp27[24], tmp27[23], tmp27[22], tmp27[21], tmp27[20], tmp27[19], tmp27[18], tmp27[17], tmp27[16], tmp27[15], tmp27[14], tmp27[13], tmp27[12], tmp27[11], tmp27[10], tmp27[9], tmp27[8], tmp27[7], tmp27[6], tmp27[5], tmp27[4], tmp27[3], tmp27[2], tmp27[1], tmp27[0]};
    assign tmp5422 = {tmp5421, const_489_0};
    assign tmp5423 = {const_490_0};
    assign tmp5424 = {tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423, tmp5423};
    assign tmp5425 = {tmp5424, const_490_0};
    assign tmp5426 = {tmp27[255]};
    assign tmp5427 = tmp5425 - tmp27;
    assign tmp5428 = {tmp5427[256]};
    assign tmp5429 = {tmp5425[255]};
    assign tmp5430 = ~tmp5429;
    assign tmp5431 = tmp5428 ^ tmp5430;
    assign tmp5432 = {tmp27[255]};
    assign tmp5433 = ~tmp5432;
    assign tmp5434 = tmp5431 ^ tmp5433;
    assign tmp5435 = {tmp5422[255]};
    assign tmp5436 = {const_491_0};
    assign tmp5437 = {tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436, tmp5436};
    assign tmp5438 = {tmp5437, const_491_0};
    assign tmp5439 = tmp5422 - tmp5438;
    assign tmp5440 = {tmp5439[256]};
    assign tmp5441 = {tmp5422[255]};
    assign tmp5442 = ~tmp5441;
    assign tmp5443 = tmp5440 ^ tmp5442;
    assign tmp5444 = {tmp5438[255]};
    assign tmp5445 = ~tmp5444;
    assign tmp5446 = tmp5443 ^ tmp5445;
    assign tmp5447 = tmp5434 & tmp5446;
    assign tmp5448 = {tmp27[255]};
    assign tmp5449 = {const_492_0};
    assign tmp5450 = {tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449, tmp5449};
    assign tmp5451 = {tmp5450, const_492_0};
    assign tmp5452 = tmp27 - tmp5451;
    assign tmp5453 = {tmp5452[256]};
    assign tmp5454 = {tmp27[255]};
    assign tmp5455 = ~tmp5454;
    assign tmp5456 = tmp5453 ^ tmp5455;
    assign tmp5457 = {tmp5451[255]};
    assign tmp5458 = ~tmp5457;
    assign tmp5459 = tmp5456 ^ tmp5458;
    assign tmp5460 = {const_493_0};
    assign tmp5461 = {tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460, tmp5460};
    assign tmp5462 = {tmp5461, const_493_0};
    assign tmp5463 = {tmp5422[255]};
    assign tmp5464 = tmp5462 - tmp5422;
    assign tmp5465 = {tmp5464[256]};
    assign tmp5466 = {tmp5462[255]};
    assign tmp5467 = ~tmp5466;
    assign tmp5468 = tmp5465 ^ tmp5467;
    assign tmp5469 = {tmp5422[255]};
    assign tmp5470 = ~tmp5469;
    assign tmp5471 = tmp5468 ^ tmp5470;
    assign tmp5472 = tmp5462 == tmp5422;
    assign tmp5473 = tmp5471 | tmp5472;
    assign tmp5474 = tmp5459 & tmp5473;
    assign tmp5475 = tmp5447 ? const_494_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp5422;
    assign tmp5476 = tmp5474 ? _ver_out_tmp_26 : tmp5475;
    assign tmp5477 = {tmp31[255]};
    assign tmp5478 = {tmp5476[255]};
    assign tmp5479 = tmp31 - tmp5476;
    assign tmp5480 = {tmp5479[256]};
    assign tmp5481 = {tmp31[255]};
    assign tmp5482 = ~tmp5481;
    assign tmp5483 = tmp5480 ^ tmp5482;
    assign tmp5484 = {tmp5476[255]};
    assign tmp5485 = ~tmp5484;
    assign tmp5486 = tmp5483 ^ tmp5485;
    assign tmp5487 = tmp5420 & tmp5486;
    assign tmp5488 = {tmp31[254], tmp31[253], tmp31[252], tmp31[251], tmp31[250], tmp31[249], tmp31[248], tmp31[247], tmp31[246], tmp31[245], tmp31[244], tmp31[243], tmp31[242], tmp31[241], tmp31[240], tmp31[239], tmp31[238], tmp31[237], tmp31[236], tmp31[235], tmp31[234], tmp31[233], tmp31[232], tmp31[231], tmp31[230], tmp31[229], tmp31[228], tmp31[227], tmp31[226], tmp31[225], tmp31[224], tmp31[223], tmp31[222], tmp31[221], tmp31[220], tmp31[219], tmp31[218], tmp31[217], tmp31[216], tmp31[215], tmp31[214], tmp31[213], tmp31[212], tmp31[211], tmp31[210], tmp31[209], tmp31[208], tmp31[207], tmp31[206], tmp31[205], tmp31[204], tmp31[203], tmp31[202], tmp31[201], tmp31[200], tmp31[199], tmp31[198], tmp31[197], tmp31[196], tmp31[195], tmp31[194], tmp31[193], tmp31[192], tmp31[191], tmp31[190], tmp31[189], tmp31[188], tmp31[187], tmp31[186], tmp31[185], tmp31[184], tmp31[183], tmp31[182], tmp31[181], tmp31[180], tmp31[179], tmp31[178], tmp31[177], tmp31[176], tmp31[175], tmp31[174], tmp31[173], tmp31[172], tmp31[171], tmp31[170], tmp31[169], tmp31[168], tmp31[167], tmp31[166], tmp31[165], tmp31[164], tmp31[163], tmp31[162], tmp31[161], tmp31[160], tmp31[159], tmp31[158], tmp31[157], tmp31[156], tmp31[155], tmp31[154], tmp31[153], tmp31[152], tmp31[151], tmp31[150], tmp31[149], tmp31[148], tmp31[147], tmp31[146], tmp31[145], tmp31[144], tmp31[143], tmp31[142], tmp31[141], tmp31[140], tmp31[139], tmp31[138], tmp31[137], tmp31[136], tmp31[135], tmp31[134], tmp31[133], tmp31[132], tmp31[131], tmp31[130], tmp31[129], tmp31[128], tmp31[127], tmp31[126], tmp31[125], tmp31[124], tmp31[123], tmp31[122], tmp31[121], tmp31[120], tmp31[119], tmp31[118], tmp31[117], tmp31[116], tmp31[115], tmp31[114], tmp31[113], tmp31[112], tmp31[111], tmp31[110], tmp31[109], tmp31[108], tmp31[107], tmp31[106], tmp31[105], tmp31[104], tmp31[103], tmp31[102], tmp31[101], tmp31[100], tmp31[99], tmp31[98], tmp31[97], tmp31[96], tmp31[95], tmp31[94], tmp31[93], tmp31[92], tmp31[91], tmp31[90], tmp31[89], tmp31[88], tmp31[87], tmp31[86], tmp31[85], tmp31[84], tmp31[83], tmp31[82], tmp31[81], tmp31[80], tmp31[79], tmp31[78], tmp31[77], tmp31[76], tmp31[75], tmp31[74], tmp31[73], tmp31[72], tmp31[71], tmp31[70], tmp31[69], tmp31[68], tmp31[67], tmp31[66], tmp31[65], tmp31[64], tmp31[63], tmp31[62], tmp31[61], tmp31[60], tmp31[59], tmp31[58], tmp31[57], tmp31[56], tmp31[55], tmp31[54], tmp31[53], tmp31[52], tmp31[51], tmp31[50], tmp31[49], tmp31[48], tmp31[47], tmp31[46], tmp31[45], tmp31[44], tmp31[43], tmp31[42], tmp31[41], tmp31[40], tmp31[39], tmp31[38], tmp31[37], tmp31[36], tmp31[35], tmp31[34], tmp31[33], tmp31[32], tmp31[31], tmp31[30], tmp31[29], tmp31[28], tmp31[27], tmp31[26], tmp31[25], tmp31[24], tmp31[23], tmp31[22], tmp31[21], tmp31[20], tmp31[19], tmp31[18], tmp31[17], tmp31[16], tmp31[15], tmp31[14], tmp31[13], tmp31[12], tmp31[11], tmp31[10], tmp31[9], tmp31[8], tmp31[7], tmp31[6], tmp31[5], tmp31[4], tmp31[3], tmp31[2], tmp31[1], tmp31[0]};
    assign tmp5489 = {tmp5488, const_496_0};
    assign tmp5490 = {const_497_0};
    assign tmp5491 = {tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490, tmp5490};
    assign tmp5492 = {tmp5491, const_497_0};
    assign tmp5493 = {tmp31[255]};
    assign tmp5494 = tmp5492 - tmp31;
    assign tmp5495 = {tmp5494[256]};
    assign tmp5496 = {tmp5492[255]};
    assign tmp5497 = ~tmp5496;
    assign tmp5498 = tmp5495 ^ tmp5497;
    assign tmp5499 = {tmp31[255]};
    assign tmp5500 = ~tmp5499;
    assign tmp5501 = tmp5498 ^ tmp5500;
    assign tmp5502 = {tmp5489[255]};
    assign tmp5503 = {const_498_0};
    assign tmp5504 = {tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503, tmp5503};
    assign tmp5505 = {tmp5504, const_498_0};
    assign tmp5506 = tmp5489 - tmp5505;
    assign tmp5507 = {tmp5506[256]};
    assign tmp5508 = {tmp5489[255]};
    assign tmp5509 = ~tmp5508;
    assign tmp5510 = tmp5507 ^ tmp5509;
    assign tmp5511 = {tmp5505[255]};
    assign tmp5512 = ~tmp5511;
    assign tmp5513 = tmp5510 ^ tmp5512;
    assign tmp5514 = tmp5501 & tmp5513;
    assign tmp5515 = {tmp31[255]};
    assign tmp5516 = {const_499_0};
    assign tmp5517 = {tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516, tmp5516};
    assign tmp5518 = {tmp5517, const_499_0};
    assign tmp5519 = tmp31 - tmp5518;
    assign tmp5520 = {tmp5519[256]};
    assign tmp5521 = {tmp31[255]};
    assign tmp5522 = ~tmp5521;
    assign tmp5523 = tmp5520 ^ tmp5522;
    assign tmp5524 = {tmp5518[255]};
    assign tmp5525 = ~tmp5524;
    assign tmp5526 = tmp5523 ^ tmp5525;
    assign tmp5527 = {const_500_0};
    assign tmp5528 = {tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527, tmp5527};
    assign tmp5529 = {tmp5528, const_500_0};
    assign tmp5530 = {tmp5489[255]};
    assign tmp5531 = tmp5529 - tmp5489;
    assign tmp5532 = {tmp5531[256]};
    assign tmp5533 = {tmp5529[255]};
    assign tmp5534 = ~tmp5533;
    assign tmp5535 = tmp5532 ^ tmp5534;
    assign tmp5536 = {tmp5489[255]};
    assign tmp5537 = ~tmp5536;
    assign tmp5538 = tmp5535 ^ tmp5537;
    assign tmp5539 = tmp5529 == tmp5489;
    assign tmp5540 = tmp5538 | tmp5539;
    assign tmp5541 = tmp5526 & tmp5540;
    assign tmp5542 = tmp5514 ? const_501_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp5489;
    assign tmp5543 = tmp5541 ? _ver_out_tmp_28 : tmp5542;
    assign tmp5544 = {tmp27[255]};
    assign tmp5545 = {tmp5543[255]};
    assign tmp5546 = tmp27 - tmp5543;
    assign tmp5547 = {tmp5546[256]};
    assign tmp5548 = {tmp27[255]};
    assign tmp5549 = ~tmp5548;
    assign tmp5550 = tmp5547 ^ tmp5549;
    assign tmp5551 = {tmp5543[255]};
    assign tmp5552 = ~tmp5551;
    assign tmp5553 = tmp5550 ^ tmp5552;
    assign tmp5554 = tmp5487 & tmp5553;
    assign tmp5555 = {tmp28[254], tmp28[253], tmp28[252], tmp28[251], tmp28[250], tmp28[249], tmp28[248], tmp28[247], tmp28[246], tmp28[245], tmp28[244], tmp28[243], tmp28[242], tmp28[241], tmp28[240], tmp28[239], tmp28[238], tmp28[237], tmp28[236], tmp28[235], tmp28[234], tmp28[233], tmp28[232], tmp28[231], tmp28[230], tmp28[229], tmp28[228], tmp28[227], tmp28[226], tmp28[225], tmp28[224], tmp28[223], tmp28[222], tmp28[221], tmp28[220], tmp28[219], tmp28[218], tmp28[217], tmp28[216], tmp28[215], tmp28[214], tmp28[213], tmp28[212], tmp28[211], tmp28[210], tmp28[209], tmp28[208], tmp28[207], tmp28[206], tmp28[205], tmp28[204], tmp28[203], tmp28[202], tmp28[201], tmp28[200], tmp28[199], tmp28[198], tmp28[197], tmp28[196], tmp28[195], tmp28[194], tmp28[193], tmp28[192], tmp28[191], tmp28[190], tmp28[189], tmp28[188], tmp28[187], tmp28[186], tmp28[185], tmp28[184], tmp28[183], tmp28[182], tmp28[181], tmp28[180], tmp28[179], tmp28[178], tmp28[177], tmp28[176], tmp28[175], tmp28[174], tmp28[173], tmp28[172], tmp28[171], tmp28[170], tmp28[169], tmp28[168], tmp28[167], tmp28[166], tmp28[165], tmp28[164], tmp28[163], tmp28[162], tmp28[161], tmp28[160], tmp28[159], tmp28[158], tmp28[157], tmp28[156], tmp28[155], tmp28[154], tmp28[153], tmp28[152], tmp28[151], tmp28[150], tmp28[149], tmp28[148], tmp28[147], tmp28[146], tmp28[145], tmp28[144], tmp28[143], tmp28[142], tmp28[141], tmp28[140], tmp28[139], tmp28[138], tmp28[137], tmp28[136], tmp28[135], tmp28[134], tmp28[133], tmp28[132], tmp28[131], tmp28[130], tmp28[129], tmp28[128], tmp28[127], tmp28[126], tmp28[125], tmp28[124], tmp28[123], tmp28[122], tmp28[121], tmp28[120], tmp28[119], tmp28[118], tmp28[117], tmp28[116], tmp28[115], tmp28[114], tmp28[113], tmp28[112], tmp28[111], tmp28[110], tmp28[109], tmp28[108], tmp28[107], tmp28[106], tmp28[105], tmp28[104], tmp28[103], tmp28[102], tmp28[101], tmp28[100], tmp28[99], tmp28[98], tmp28[97], tmp28[96], tmp28[95], tmp28[94], tmp28[93], tmp28[92], tmp28[91], tmp28[90], tmp28[89], tmp28[88], tmp28[87], tmp28[86], tmp28[85], tmp28[84], tmp28[83], tmp28[82], tmp28[81], tmp28[80], tmp28[79], tmp28[78], tmp28[77], tmp28[76], tmp28[75], tmp28[74], tmp28[73], tmp28[72], tmp28[71], tmp28[70], tmp28[69], tmp28[68], tmp28[67], tmp28[66], tmp28[65], tmp28[64], tmp28[63], tmp28[62], tmp28[61], tmp28[60], tmp28[59], tmp28[58], tmp28[57], tmp28[56], tmp28[55], tmp28[54], tmp28[53], tmp28[52], tmp28[51], tmp28[50], tmp28[49], tmp28[48], tmp28[47], tmp28[46], tmp28[45], tmp28[44], tmp28[43], tmp28[42], tmp28[41], tmp28[40], tmp28[39], tmp28[38], tmp28[37], tmp28[36], tmp28[35], tmp28[34], tmp28[33], tmp28[32], tmp28[31], tmp28[30], tmp28[29], tmp28[28], tmp28[27], tmp28[26], tmp28[25], tmp28[24], tmp28[23], tmp28[22], tmp28[21], tmp28[20], tmp28[19], tmp28[18], tmp28[17], tmp28[16], tmp28[15], tmp28[14], tmp28[13], tmp28[12], tmp28[11], tmp28[10], tmp28[9], tmp28[8], tmp28[7], tmp28[6], tmp28[5], tmp28[4], tmp28[3], tmp28[2], tmp28[1], tmp28[0]};
    assign tmp5556 = {tmp5555, const_503_0};
    assign tmp5557 = {const_504_0};
    assign tmp5558 = {tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557, tmp5557};
    assign tmp5559 = {tmp5558, const_504_0};
    assign tmp5560 = {tmp28[255]};
    assign tmp5561 = tmp5559 - tmp28;
    assign tmp5562 = {tmp5561[256]};
    assign tmp5563 = {tmp5559[255]};
    assign tmp5564 = ~tmp5563;
    assign tmp5565 = tmp5562 ^ tmp5564;
    assign tmp5566 = {tmp28[255]};
    assign tmp5567 = ~tmp5566;
    assign tmp5568 = tmp5565 ^ tmp5567;
    assign tmp5569 = {tmp5556[255]};
    assign tmp5570 = {const_505_0};
    assign tmp5571 = {tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570, tmp5570};
    assign tmp5572 = {tmp5571, const_505_0};
    assign tmp5573 = tmp5556 - tmp5572;
    assign tmp5574 = {tmp5573[256]};
    assign tmp5575 = {tmp5556[255]};
    assign tmp5576 = ~tmp5575;
    assign tmp5577 = tmp5574 ^ tmp5576;
    assign tmp5578 = {tmp5572[255]};
    assign tmp5579 = ~tmp5578;
    assign tmp5580 = tmp5577 ^ tmp5579;
    assign tmp5581 = tmp5568 & tmp5580;
    assign tmp5582 = {tmp28[255]};
    assign tmp5583 = {const_506_0};
    assign tmp5584 = {tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583, tmp5583};
    assign tmp5585 = {tmp5584, const_506_0};
    assign tmp5586 = tmp28 - tmp5585;
    assign tmp5587 = {tmp5586[256]};
    assign tmp5588 = {tmp28[255]};
    assign tmp5589 = ~tmp5588;
    assign tmp5590 = tmp5587 ^ tmp5589;
    assign tmp5591 = {tmp5585[255]};
    assign tmp5592 = ~tmp5591;
    assign tmp5593 = tmp5590 ^ tmp5592;
    assign tmp5594 = {const_507_0};
    assign tmp5595 = {tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594, tmp5594};
    assign tmp5596 = {tmp5595, const_507_0};
    assign tmp5597 = {tmp5556[255]};
    assign tmp5598 = tmp5596 - tmp5556;
    assign tmp5599 = {tmp5598[256]};
    assign tmp5600 = {tmp5596[255]};
    assign tmp5601 = ~tmp5600;
    assign tmp5602 = tmp5599 ^ tmp5601;
    assign tmp5603 = {tmp5556[255]};
    assign tmp5604 = ~tmp5603;
    assign tmp5605 = tmp5602 ^ tmp5604;
    assign tmp5606 = tmp5596 == tmp5556;
    assign tmp5607 = tmp5605 | tmp5606;
    assign tmp5608 = tmp5593 & tmp5607;
    assign tmp5609 = tmp5581 ? const_508_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp5556;
    assign tmp5610 = tmp5608 ? _ver_out_tmp_31 : tmp5609;
    assign tmp5611 = {tmp32[255]};
    assign tmp5612 = {tmp5610[255]};
    assign tmp5613 = tmp32 - tmp5610;
    assign tmp5614 = {tmp5613[256]};
    assign tmp5615 = {tmp32[255]};
    assign tmp5616 = ~tmp5615;
    assign tmp5617 = tmp5614 ^ tmp5616;
    assign tmp5618 = {tmp5610[255]};
    assign tmp5619 = ~tmp5618;
    assign tmp5620 = tmp5617 ^ tmp5619;
    assign tmp5621 = tmp5554 & tmp5620;
    assign tmp5622 = {tmp32[254], tmp32[253], tmp32[252], tmp32[251], tmp32[250], tmp32[249], tmp32[248], tmp32[247], tmp32[246], tmp32[245], tmp32[244], tmp32[243], tmp32[242], tmp32[241], tmp32[240], tmp32[239], tmp32[238], tmp32[237], tmp32[236], tmp32[235], tmp32[234], tmp32[233], tmp32[232], tmp32[231], tmp32[230], tmp32[229], tmp32[228], tmp32[227], tmp32[226], tmp32[225], tmp32[224], tmp32[223], tmp32[222], tmp32[221], tmp32[220], tmp32[219], tmp32[218], tmp32[217], tmp32[216], tmp32[215], tmp32[214], tmp32[213], tmp32[212], tmp32[211], tmp32[210], tmp32[209], tmp32[208], tmp32[207], tmp32[206], tmp32[205], tmp32[204], tmp32[203], tmp32[202], tmp32[201], tmp32[200], tmp32[199], tmp32[198], tmp32[197], tmp32[196], tmp32[195], tmp32[194], tmp32[193], tmp32[192], tmp32[191], tmp32[190], tmp32[189], tmp32[188], tmp32[187], tmp32[186], tmp32[185], tmp32[184], tmp32[183], tmp32[182], tmp32[181], tmp32[180], tmp32[179], tmp32[178], tmp32[177], tmp32[176], tmp32[175], tmp32[174], tmp32[173], tmp32[172], tmp32[171], tmp32[170], tmp32[169], tmp32[168], tmp32[167], tmp32[166], tmp32[165], tmp32[164], tmp32[163], tmp32[162], tmp32[161], tmp32[160], tmp32[159], tmp32[158], tmp32[157], tmp32[156], tmp32[155], tmp32[154], tmp32[153], tmp32[152], tmp32[151], tmp32[150], tmp32[149], tmp32[148], tmp32[147], tmp32[146], tmp32[145], tmp32[144], tmp32[143], tmp32[142], tmp32[141], tmp32[140], tmp32[139], tmp32[138], tmp32[137], tmp32[136], tmp32[135], tmp32[134], tmp32[133], tmp32[132], tmp32[131], tmp32[130], tmp32[129], tmp32[128], tmp32[127], tmp32[126], tmp32[125], tmp32[124], tmp32[123], tmp32[122], tmp32[121], tmp32[120], tmp32[119], tmp32[118], tmp32[117], tmp32[116], tmp32[115], tmp32[114], tmp32[113], tmp32[112], tmp32[111], tmp32[110], tmp32[109], tmp32[108], tmp32[107], tmp32[106], tmp32[105], tmp32[104], tmp32[103], tmp32[102], tmp32[101], tmp32[100], tmp32[99], tmp32[98], tmp32[97], tmp32[96], tmp32[95], tmp32[94], tmp32[93], tmp32[92], tmp32[91], tmp32[90], tmp32[89], tmp32[88], tmp32[87], tmp32[86], tmp32[85], tmp32[84], tmp32[83], tmp32[82], tmp32[81], tmp32[80], tmp32[79], tmp32[78], tmp32[77], tmp32[76], tmp32[75], tmp32[74], tmp32[73], tmp32[72], tmp32[71], tmp32[70], tmp32[69], tmp32[68], tmp32[67], tmp32[66], tmp32[65], tmp32[64], tmp32[63], tmp32[62], tmp32[61], tmp32[60], tmp32[59], tmp32[58], tmp32[57], tmp32[56], tmp32[55], tmp32[54], tmp32[53], tmp32[52], tmp32[51], tmp32[50], tmp32[49], tmp32[48], tmp32[47], tmp32[46], tmp32[45], tmp32[44], tmp32[43], tmp32[42], tmp32[41], tmp32[40], tmp32[39], tmp32[38], tmp32[37], tmp32[36], tmp32[35], tmp32[34], tmp32[33], tmp32[32], tmp32[31], tmp32[30], tmp32[29], tmp32[28], tmp32[27], tmp32[26], tmp32[25], tmp32[24], tmp32[23], tmp32[22], tmp32[21], tmp32[20], tmp32[19], tmp32[18], tmp32[17], tmp32[16], tmp32[15], tmp32[14], tmp32[13], tmp32[12], tmp32[11], tmp32[10], tmp32[9], tmp32[8], tmp32[7], tmp32[6], tmp32[5], tmp32[4], tmp32[3], tmp32[2], tmp32[1], tmp32[0]};
    assign tmp5623 = {tmp5622, const_510_0};
    assign tmp5624 = {const_511_0};
    assign tmp5625 = {tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624, tmp5624};
    assign tmp5626 = {tmp5625, const_511_0};
    assign tmp5627 = {tmp32[255]};
    assign tmp5628 = tmp5626 - tmp32;
    assign tmp5629 = {tmp5628[256]};
    assign tmp5630 = {tmp5626[255]};
    assign tmp5631 = ~tmp5630;
    assign tmp5632 = tmp5629 ^ tmp5631;
    assign tmp5633 = {tmp32[255]};
    assign tmp5634 = ~tmp5633;
    assign tmp5635 = tmp5632 ^ tmp5634;
    assign tmp5636 = {tmp5623[255]};
    assign tmp5637 = {const_512_0};
    assign tmp5638 = {tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637, tmp5637};
    assign tmp5639 = {tmp5638, const_512_0};
    assign tmp5640 = tmp5623 - tmp5639;
    assign tmp5641 = {tmp5640[256]};
    assign tmp5642 = {tmp5623[255]};
    assign tmp5643 = ~tmp5642;
    assign tmp5644 = tmp5641 ^ tmp5643;
    assign tmp5645 = {tmp5639[255]};
    assign tmp5646 = ~tmp5645;
    assign tmp5647 = tmp5644 ^ tmp5646;
    assign tmp5648 = tmp5635 & tmp5647;
    assign tmp5649 = {tmp32[255]};
    assign tmp5650 = {const_513_0};
    assign tmp5651 = {tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650, tmp5650};
    assign tmp5652 = {tmp5651, const_513_0};
    assign tmp5653 = tmp32 - tmp5652;
    assign tmp5654 = {tmp5653[256]};
    assign tmp5655 = {tmp32[255]};
    assign tmp5656 = ~tmp5655;
    assign tmp5657 = tmp5654 ^ tmp5656;
    assign tmp5658 = {tmp5652[255]};
    assign tmp5659 = ~tmp5658;
    assign tmp5660 = tmp5657 ^ tmp5659;
    assign tmp5661 = {const_514_0};
    assign tmp5662 = {tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661, tmp5661};
    assign tmp5663 = {tmp5662, const_514_0};
    assign tmp5664 = {tmp5623[255]};
    assign tmp5665 = tmp5663 - tmp5623;
    assign tmp5666 = {tmp5665[256]};
    assign tmp5667 = {tmp5663[255]};
    assign tmp5668 = ~tmp5667;
    assign tmp5669 = tmp5666 ^ tmp5668;
    assign tmp5670 = {tmp5623[255]};
    assign tmp5671 = ~tmp5670;
    assign tmp5672 = tmp5669 ^ tmp5671;
    assign tmp5673 = tmp5663 == tmp5623;
    assign tmp5674 = tmp5672 | tmp5673;
    assign tmp5675 = tmp5660 & tmp5674;
    assign tmp5676 = tmp5648 ? const_515_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp5623;
    assign tmp5677 = tmp5675 ? _ver_out_tmp_35 : tmp5676;
    assign tmp5678 = {tmp28[255]};
    assign tmp5679 = {tmp5677[255]};
    assign tmp5680 = tmp28 - tmp5677;
    assign tmp5681 = {tmp5680[256]};
    assign tmp5682 = {tmp28[255]};
    assign tmp5683 = ~tmp5682;
    assign tmp5684 = tmp5681 ^ tmp5683;
    assign tmp5685 = {tmp5677[255]};
    assign tmp5686 = ~tmp5685;
    assign tmp5687 = tmp5684 ^ tmp5686;
    assign tmp5688 = tmp5621 & tmp5687;
    assign tmp5689 = ~tmp35;
    assign tmp5690 = ~tmp36;
    assign tmp5691 = tmp5689 & tmp5690;
    assign tmp5692 = ~tmp57;
    assign tmp5693 = tmp5691 & tmp5692;
    assign tmp5694 = ~tmp1034;
    assign tmp5695 = tmp5693 & tmp5694;
    assign tmp5696 = tmp5695 & tmp2071;
    assign tmp5697 = ~tmp2583;
    assign tmp5698 = tmp5696 & tmp5697;
    assign tmp5699 = tmp5698 & tmp23;
    assign tmp5700 = ~tmp2627;
    assign tmp5701 = tmp5699 & tmp5700;
    assign tmp5702 = ~tmp2798;
    assign tmp5703 = tmp5701 & tmp5702;
    assign tmp5704 = ~tmp3425;
    assign tmp5705 = tmp5703 & tmp5704;
    assign tmp5706 = ~tmp4020;
    assign tmp5707 = tmp5705 & tmp5706;
    assign tmp5708 = tmp5707 & cfg_speculative_egest;
    assign tmp5709 = ~tmp4511;
    assign tmp5710 = tmp5708 & tmp5709;
    assign tmp5711 = tmp5710 & tmp5688;
    assign tmp5712 = ~tmp35;
    assign tmp5713 = ~tmp36;
    assign tmp5714 = tmp5712 & tmp5713;
    assign tmp5715 = ~tmp57;
    assign tmp5716 = tmp5714 & tmp5715;
    assign tmp5717 = ~tmp1034;
    assign tmp5718 = tmp5716 & tmp5717;
    assign tmp5719 = tmp5718 & tmp2071;
    assign tmp5720 = ~tmp2583;
    assign tmp5721 = tmp5719 & tmp5720;
    assign tmp5722 = tmp5721 & tmp23;
    assign tmp5723 = ~tmp2627;
    assign tmp5724 = tmp5722 & tmp5723;
    assign tmp5725 = ~tmp2798;
    assign tmp5726 = tmp5724 & tmp5725;
    assign tmp5727 = ~tmp3425;
    assign tmp5728 = tmp5726 & tmp5727;
    assign tmp5729 = ~tmp4020;
    assign tmp5730 = tmp5728 & tmp5729;
    assign tmp5731 = tmp5730 & cfg_speculative_egest;
    assign tmp5732 = ~tmp4511;
    assign tmp5733 = tmp5731 & tmp5732;
    assign tmp5734 = tmp5733 & tmp5688;
    assign tmp5735 = ~tmp35;
    assign tmp5736 = ~tmp36;
    assign tmp5737 = tmp5735 & tmp5736;
    assign tmp5738 = ~tmp57;
    assign tmp5739 = tmp5737 & tmp5738;
    assign tmp5740 = ~tmp1034;
    assign tmp5741 = tmp5739 & tmp5740;
    assign tmp5742 = tmp5741 & tmp2071;
    assign tmp5743 = ~tmp2583;
    assign tmp5744 = tmp5742 & tmp5743;
    assign tmp5745 = tmp5744 & tmp23;
    assign tmp5746 = ~tmp2627;
    assign tmp5747 = tmp5745 & tmp5746;
    assign tmp5748 = ~tmp2798;
    assign tmp5749 = tmp5747 & tmp5748;
    assign tmp5750 = ~tmp3425;
    assign tmp5751 = tmp5749 & tmp5750;
    assign tmp5752 = ~tmp4020;
    assign tmp5753 = tmp5751 & tmp5752;
    assign tmp5754 = tmp5753 & cfg_speculative_egest;
    assign tmp5755 = ~tmp4511;
    assign tmp5756 = tmp5754 & tmp5755;
    assign tmp5757 = tmp5756 & tmp5688;
    assign tmp5758 = _ver_out_tmp_37 == tmp29;
    assign tmp5759 = {const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0, const_521_0};
    assign tmp5760 = {tmp5759, const_520_0};
    assign tmp5761 = tmp5760 - tmp29;
    assign tmp5762 = {const_523_0, const_523_0};
    assign tmp5763 = {tmp5762, const_522_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp5764 = tmp5758 ? tmp5763 : tmp5761;
    assign tmp5765 = {tmp25[255]};
    assign tmp5766 = {tmp5765, tmp5765};
    assign tmp5767 = {tmp5766, tmp25};
    assign tmp5768 = {tmp5764[256]};
    assign tmp5769 = {tmp5768};
    assign tmp5770 = {tmp5769, tmp5764};
    assign tmp5771 = tmp5767 + tmp5770;
    assign tmp5772 = {tmp5771[257], tmp5771[256], tmp5771[255], tmp5771[254], tmp5771[253], tmp5771[252], tmp5771[251], tmp5771[250], tmp5771[249], tmp5771[248], tmp5771[247], tmp5771[246], tmp5771[245], tmp5771[244], tmp5771[243], tmp5771[242], tmp5771[241], tmp5771[240], tmp5771[239], tmp5771[238], tmp5771[237], tmp5771[236], tmp5771[235], tmp5771[234], tmp5771[233], tmp5771[232], tmp5771[231], tmp5771[230], tmp5771[229], tmp5771[228], tmp5771[227], tmp5771[226], tmp5771[225], tmp5771[224], tmp5771[223], tmp5771[222], tmp5771[221], tmp5771[220], tmp5771[219], tmp5771[218], tmp5771[217], tmp5771[216], tmp5771[215], tmp5771[214], tmp5771[213], tmp5771[212], tmp5771[211], tmp5771[210], tmp5771[209], tmp5771[208], tmp5771[207], tmp5771[206], tmp5771[205], tmp5771[204], tmp5771[203], tmp5771[202], tmp5771[201], tmp5771[200], tmp5771[199], tmp5771[198], tmp5771[197], tmp5771[196], tmp5771[195], tmp5771[194], tmp5771[193], tmp5771[192], tmp5771[191], tmp5771[190], tmp5771[189], tmp5771[188], tmp5771[187], tmp5771[186], tmp5771[185], tmp5771[184], tmp5771[183], tmp5771[182], tmp5771[181], tmp5771[180], tmp5771[179], tmp5771[178], tmp5771[177], tmp5771[176], tmp5771[175], tmp5771[174], tmp5771[173], tmp5771[172], tmp5771[171], tmp5771[170], tmp5771[169], tmp5771[168], tmp5771[167], tmp5771[166], tmp5771[165], tmp5771[164], tmp5771[163], tmp5771[162], tmp5771[161], tmp5771[160], tmp5771[159], tmp5771[158], tmp5771[157], tmp5771[156], tmp5771[155], tmp5771[154], tmp5771[153], tmp5771[152], tmp5771[151], tmp5771[150], tmp5771[149], tmp5771[148], tmp5771[147], tmp5771[146], tmp5771[145], tmp5771[144], tmp5771[143], tmp5771[142], tmp5771[141], tmp5771[140], tmp5771[139], tmp5771[138], tmp5771[137], tmp5771[136], tmp5771[135], tmp5771[134], tmp5771[133], tmp5771[132], tmp5771[131], tmp5771[130], tmp5771[129], tmp5771[128], tmp5771[127], tmp5771[126], tmp5771[125], tmp5771[124], tmp5771[123], tmp5771[122], tmp5771[121], tmp5771[120], tmp5771[119], tmp5771[118], tmp5771[117], tmp5771[116], tmp5771[115], tmp5771[114], tmp5771[113], tmp5771[112], tmp5771[111], tmp5771[110], tmp5771[109], tmp5771[108], tmp5771[107], tmp5771[106], tmp5771[105], tmp5771[104], tmp5771[103], tmp5771[102], tmp5771[101], tmp5771[100], tmp5771[99], tmp5771[98], tmp5771[97], tmp5771[96], tmp5771[95], tmp5771[94], tmp5771[93], tmp5771[92], tmp5771[91], tmp5771[90], tmp5771[89], tmp5771[88], tmp5771[87], tmp5771[86], tmp5771[85], tmp5771[84], tmp5771[83], tmp5771[82], tmp5771[81], tmp5771[80], tmp5771[79], tmp5771[78], tmp5771[77], tmp5771[76], tmp5771[75], tmp5771[74], tmp5771[73], tmp5771[72], tmp5771[71], tmp5771[70], tmp5771[69], tmp5771[68], tmp5771[67], tmp5771[66], tmp5771[65], tmp5771[64], tmp5771[63], tmp5771[62], tmp5771[61], tmp5771[60], tmp5771[59], tmp5771[58], tmp5771[57], tmp5771[56], tmp5771[55], tmp5771[54], tmp5771[53], tmp5771[52], tmp5771[51], tmp5771[50], tmp5771[49], tmp5771[48], tmp5771[47], tmp5771[46], tmp5771[45], tmp5771[44], tmp5771[43], tmp5771[42], tmp5771[41], tmp5771[40], tmp5771[39], tmp5771[38], tmp5771[37], tmp5771[36], tmp5771[35], tmp5771[34], tmp5771[33], tmp5771[32], tmp5771[31], tmp5771[30], tmp5771[29], tmp5771[28], tmp5771[27], tmp5771[26], tmp5771[25], tmp5771[24], tmp5771[23], tmp5771[22], tmp5771[21], tmp5771[20], tmp5771[19], tmp5771[18], tmp5771[17], tmp5771[16], tmp5771[15], tmp5771[14], tmp5771[13], tmp5771[12], tmp5771[11], tmp5771[10], tmp5771[9], tmp5771[8], tmp5771[7], tmp5771[6], tmp5771[5], tmp5771[4], tmp5771[3], tmp5771[2], tmp5771[1], tmp5771[0]};
    assign tmp5773 = {tmp5772[255], tmp5772[254], tmp5772[253], tmp5772[252], tmp5772[251], tmp5772[250], tmp5772[249], tmp5772[248], tmp5772[247], tmp5772[246], tmp5772[245], tmp5772[244], tmp5772[243], tmp5772[242], tmp5772[241], tmp5772[240], tmp5772[239], tmp5772[238], tmp5772[237], tmp5772[236], tmp5772[235], tmp5772[234], tmp5772[233], tmp5772[232], tmp5772[231], tmp5772[230], tmp5772[229], tmp5772[228], tmp5772[227], tmp5772[226], tmp5772[225], tmp5772[224], tmp5772[223], tmp5772[222], tmp5772[221], tmp5772[220], tmp5772[219], tmp5772[218], tmp5772[217], tmp5772[216], tmp5772[215], tmp5772[214], tmp5772[213], tmp5772[212], tmp5772[211], tmp5772[210], tmp5772[209], tmp5772[208], tmp5772[207], tmp5772[206], tmp5772[205], tmp5772[204], tmp5772[203], tmp5772[202], tmp5772[201], tmp5772[200], tmp5772[199], tmp5772[198], tmp5772[197], tmp5772[196], tmp5772[195], tmp5772[194], tmp5772[193], tmp5772[192], tmp5772[191], tmp5772[190], tmp5772[189], tmp5772[188], tmp5772[187], tmp5772[186], tmp5772[185], tmp5772[184], tmp5772[183], tmp5772[182], tmp5772[181], tmp5772[180], tmp5772[179], tmp5772[178], tmp5772[177], tmp5772[176], tmp5772[175], tmp5772[174], tmp5772[173], tmp5772[172], tmp5772[171], tmp5772[170], tmp5772[169], tmp5772[168], tmp5772[167], tmp5772[166], tmp5772[165], tmp5772[164], tmp5772[163], tmp5772[162], tmp5772[161], tmp5772[160], tmp5772[159], tmp5772[158], tmp5772[157], tmp5772[156], tmp5772[155], tmp5772[154], tmp5772[153], tmp5772[152], tmp5772[151], tmp5772[150], tmp5772[149], tmp5772[148], tmp5772[147], tmp5772[146], tmp5772[145], tmp5772[144], tmp5772[143], tmp5772[142], tmp5772[141], tmp5772[140], tmp5772[139], tmp5772[138], tmp5772[137], tmp5772[136], tmp5772[135], tmp5772[134], tmp5772[133], tmp5772[132], tmp5772[131], tmp5772[130], tmp5772[129], tmp5772[128], tmp5772[127], tmp5772[126], tmp5772[125], tmp5772[124], tmp5772[123], tmp5772[122], tmp5772[121], tmp5772[120], tmp5772[119], tmp5772[118], tmp5772[117], tmp5772[116], tmp5772[115], tmp5772[114], tmp5772[113], tmp5772[112], tmp5772[111], tmp5772[110], tmp5772[109], tmp5772[108], tmp5772[107], tmp5772[106], tmp5772[105], tmp5772[104], tmp5772[103], tmp5772[102], tmp5772[101], tmp5772[100], tmp5772[99], tmp5772[98], tmp5772[97], tmp5772[96], tmp5772[95], tmp5772[94], tmp5772[93], tmp5772[92], tmp5772[91], tmp5772[90], tmp5772[89], tmp5772[88], tmp5772[87], tmp5772[86], tmp5772[85], tmp5772[84], tmp5772[83], tmp5772[82], tmp5772[81], tmp5772[80], tmp5772[79], tmp5772[78], tmp5772[77], tmp5772[76], tmp5772[75], tmp5772[74], tmp5772[73], tmp5772[72], tmp5772[71], tmp5772[70], tmp5772[69], tmp5772[68], tmp5772[67], tmp5772[66], tmp5772[65], tmp5772[64], tmp5772[63], tmp5772[62], tmp5772[61], tmp5772[60], tmp5772[59], tmp5772[58], tmp5772[57], tmp5772[56], tmp5772[55], tmp5772[54], tmp5772[53], tmp5772[52], tmp5772[51], tmp5772[50], tmp5772[49], tmp5772[48], tmp5772[47], tmp5772[46], tmp5772[45], tmp5772[44], tmp5772[43], tmp5772[42], tmp5772[41], tmp5772[40], tmp5772[39], tmp5772[38], tmp5772[37], tmp5772[36], tmp5772[35], tmp5772[34], tmp5772[33], tmp5772[32], tmp5772[31], tmp5772[30], tmp5772[29], tmp5772[28], tmp5772[27], tmp5772[26], tmp5772[25], tmp5772[24], tmp5772[23], tmp5772[22], tmp5772[21], tmp5772[20], tmp5772[19], tmp5772[18], tmp5772[17], tmp5772[16], tmp5772[15], tmp5772[14], tmp5772[13], tmp5772[12], tmp5772[11], tmp5772[10], tmp5772[9], tmp5772[8], tmp5772[7], tmp5772[6], tmp5772[5], tmp5772[4], tmp5772[3], tmp5772[2], tmp5772[1], tmp5772[0]};
    assign tmp5774 = {const_524_0};
    assign tmp5775 = {tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774, tmp5774};
    assign tmp5776 = {tmp5775, const_524_0};
    assign tmp5777 = {tmp25[255]};
    assign tmp5778 = tmp5776 - tmp25;
    assign tmp5779 = {tmp5778[256]};
    assign tmp5780 = {tmp5776[255]};
    assign tmp5781 = ~tmp5780;
    assign tmp5782 = tmp5779 ^ tmp5781;
    assign tmp5783 = {tmp25[255]};
    assign tmp5784 = ~tmp5783;
    assign tmp5785 = tmp5782 ^ tmp5784;
    assign tmp5786 = {const_525_0};
    assign tmp5787 = {tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786, tmp5786};
    assign tmp5788 = {tmp5787, const_525_0};
    assign tmp5789 = {tmp5764[256]};
    assign tmp5790 = tmp5788 - tmp5764;
    assign tmp5791 = {tmp5790[257]};
    assign tmp5792 = {tmp5788[256]};
    assign tmp5793 = ~tmp5792;
    assign tmp5794 = tmp5791 ^ tmp5793;
    assign tmp5795 = {tmp5764[256]};
    assign tmp5796 = ~tmp5795;
    assign tmp5797 = tmp5794 ^ tmp5796;
    assign tmp5798 = tmp5785 & tmp5797;
    assign tmp5799 = {tmp5773[255]};
    assign tmp5800 = {const_526_0};
    assign tmp5801 = {tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800, tmp5800};
    assign tmp5802 = {tmp5801, const_526_0};
    assign tmp5803 = tmp5773 - tmp5802;
    assign tmp5804 = {tmp5803[256]};
    assign tmp5805 = {tmp5773[255]};
    assign tmp5806 = ~tmp5805;
    assign tmp5807 = tmp5804 ^ tmp5806;
    assign tmp5808 = {tmp5802[255]};
    assign tmp5809 = ~tmp5808;
    assign tmp5810 = tmp5807 ^ tmp5809;
    assign tmp5811 = tmp5773 == tmp5802;
    assign tmp5812 = tmp5810 | tmp5811;
    assign tmp5813 = tmp5798 & tmp5812;
    assign tmp5814 = {tmp25[255]};
    assign tmp5815 = {const_527_0};
    assign tmp5816 = {tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815, tmp5815};
    assign tmp5817 = {tmp5816, const_527_0};
    assign tmp5818 = tmp25 - tmp5817;
    assign tmp5819 = {tmp5818[256]};
    assign tmp5820 = {tmp25[255]};
    assign tmp5821 = ~tmp5820;
    assign tmp5822 = tmp5819 ^ tmp5821;
    assign tmp5823 = {tmp5817[255]};
    assign tmp5824 = ~tmp5823;
    assign tmp5825 = tmp5822 ^ tmp5824;
    assign tmp5826 = {tmp5764[256]};
    assign tmp5827 = {const_528_0};
    assign tmp5828 = {tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827, tmp5827};
    assign tmp5829 = {tmp5828, const_528_0};
    assign tmp5830 = tmp5764 - tmp5829;
    assign tmp5831 = {tmp5830[257]};
    assign tmp5832 = {tmp5764[256]};
    assign tmp5833 = ~tmp5832;
    assign tmp5834 = tmp5831 ^ tmp5833;
    assign tmp5835 = {tmp5829[256]};
    assign tmp5836 = ~tmp5835;
    assign tmp5837 = tmp5834 ^ tmp5836;
    assign tmp5838 = tmp5825 & tmp5837;
    assign tmp5839 = {const_529_0};
    assign tmp5840 = {tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839, tmp5839};
    assign tmp5841 = {tmp5840, const_529_0};
    assign tmp5842 = {tmp5773[255]};
    assign tmp5843 = tmp5841 - tmp5773;
    assign tmp5844 = {tmp5843[256]};
    assign tmp5845 = {tmp5841[255]};
    assign tmp5846 = ~tmp5845;
    assign tmp5847 = tmp5844 ^ tmp5846;
    assign tmp5848 = {tmp5773[255]};
    assign tmp5849 = ~tmp5848;
    assign tmp5850 = tmp5847 ^ tmp5849;
    assign tmp5851 = tmp5841 == tmp5773;
    assign tmp5852 = tmp5850 | tmp5851;
    assign tmp5853 = tmp5838 & tmp5852;
    assign tmp5854 = tmp5813 ? const_530_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp5773;
    assign tmp5855 = tmp5853 ? _ver_out_tmp_42 : tmp5854;
    assign tmp5856 = ~tmp35;
    assign tmp5857 = ~tmp36;
    assign tmp5858 = tmp5856 & tmp5857;
    assign tmp5859 = ~tmp57;
    assign tmp5860 = tmp5858 & tmp5859;
    assign tmp5861 = ~tmp1034;
    assign tmp5862 = tmp5860 & tmp5861;
    assign tmp5863 = tmp5862 & tmp2071;
    assign tmp5864 = ~tmp2583;
    assign tmp5865 = tmp5863 & tmp5864;
    assign tmp5866 = tmp5865 & tmp23;
    assign tmp5867 = ~tmp2627;
    assign tmp5868 = tmp5866 & tmp5867;
    assign tmp5869 = ~tmp2798;
    assign tmp5870 = tmp5868 & tmp5869;
    assign tmp5871 = ~tmp3425;
    assign tmp5872 = tmp5870 & tmp5871;
    assign tmp5873 = ~tmp4020;
    assign tmp5874 = tmp5872 & tmp5873;
    assign tmp5875 = tmp5874 & cfg_speculative_egest;
    assign tmp5876 = ~tmp4511;
    assign tmp5877 = tmp5875 & tmp5876;
    assign tmp5878 = tmp5877 & tmp5688;
    assign tmp5879 = ~tmp35;
    assign tmp5880 = ~tmp36;
    assign tmp5881 = tmp5879 & tmp5880;
    assign tmp5882 = ~tmp57;
    assign tmp5883 = tmp5881 & tmp5882;
    assign tmp5884 = ~tmp1034;
    assign tmp5885 = tmp5883 & tmp5884;
    assign tmp5886 = tmp5885 & tmp2071;
    assign tmp5887 = ~tmp2583;
    assign tmp5888 = tmp5886 & tmp5887;
    assign tmp5889 = tmp5888 & tmp23;
    assign tmp5890 = ~tmp2627;
    assign tmp5891 = tmp5889 & tmp5890;
    assign tmp5892 = ~tmp2798;
    assign tmp5893 = tmp5891 & tmp5892;
    assign tmp5894 = ~tmp3425;
    assign tmp5895 = tmp5893 & tmp5894;
    assign tmp5896 = ~tmp4020;
    assign tmp5897 = tmp5895 & tmp5896;
    assign tmp5898 = tmp5897 & cfg_speculative_egest;
    assign tmp5899 = ~tmp4511;
    assign tmp5900 = tmp5898 & tmp5899;
    assign tmp5901 = tmp5900 & tmp5688;
    assign tmp5902 = _ver_out_tmp_44 == tmp30;
    assign tmp5903 = {const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0, const_534_0};
    assign tmp5904 = {tmp5903, const_533_0};
    assign tmp5905 = tmp5904 - tmp30;
    assign tmp5906 = {const_536_0, const_536_0};
    assign tmp5907 = {tmp5906, const_535_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp5908 = tmp5902 ? tmp5907 : tmp5905;
    assign tmp5909 = {tmp26[255]};
    assign tmp5910 = {tmp5909, tmp5909};
    assign tmp5911 = {tmp5910, tmp26};
    assign tmp5912 = {tmp5908[256]};
    assign tmp5913 = {tmp5912};
    assign tmp5914 = {tmp5913, tmp5908};
    assign tmp5915 = tmp5911 + tmp5914;
    assign tmp5916 = {tmp5915[257], tmp5915[256], tmp5915[255], tmp5915[254], tmp5915[253], tmp5915[252], tmp5915[251], tmp5915[250], tmp5915[249], tmp5915[248], tmp5915[247], tmp5915[246], tmp5915[245], tmp5915[244], tmp5915[243], tmp5915[242], tmp5915[241], tmp5915[240], tmp5915[239], tmp5915[238], tmp5915[237], tmp5915[236], tmp5915[235], tmp5915[234], tmp5915[233], tmp5915[232], tmp5915[231], tmp5915[230], tmp5915[229], tmp5915[228], tmp5915[227], tmp5915[226], tmp5915[225], tmp5915[224], tmp5915[223], tmp5915[222], tmp5915[221], tmp5915[220], tmp5915[219], tmp5915[218], tmp5915[217], tmp5915[216], tmp5915[215], tmp5915[214], tmp5915[213], tmp5915[212], tmp5915[211], tmp5915[210], tmp5915[209], tmp5915[208], tmp5915[207], tmp5915[206], tmp5915[205], tmp5915[204], tmp5915[203], tmp5915[202], tmp5915[201], tmp5915[200], tmp5915[199], tmp5915[198], tmp5915[197], tmp5915[196], tmp5915[195], tmp5915[194], tmp5915[193], tmp5915[192], tmp5915[191], tmp5915[190], tmp5915[189], tmp5915[188], tmp5915[187], tmp5915[186], tmp5915[185], tmp5915[184], tmp5915[183], tmp5915[182], tmp5915[181], tmp5915[180], tmp5915[179], tmp5915[178], tmp5915[177], tmp5915[176], tmp5915[175], tmp5915[174], tmp5915[173], tmp5915[172], tmp5915[171], tmp5915[170], tmp5915[169], tmp5915[168], tmp5915[167], tmp5915[166], tmp5915[165], tmp5915[164], tmp5915[163], tmp5915[162], tmp5915[161], tmp5915[160], tmp5915[159], tmp5915[158], tmp5915[157], tmp5915[156], tmp5915[155], tmp5915[154], tmp5915[153], tmp5915[152], tmp5915[151], tmp5915[150], tmp5915[149], tmp5915[148], tmp5915[147], tmp5915[146], tmp5915[145], tmp5915[144], tmp5915[143], tmp5915[142], tmp5915[141], tmp5915[140], tmp5915[139], tmp5915[138], tmp5915[137], tmp5915[136], tmp5915[135], tmp5915[134], tmp5915[133], tmp5915[132], tmp5915[131], tmp5915[130], tmp5915[129], tmp5915[128], tmp5915[127], tmp5915[126], tmp5915[125], tmp5915[124], tmp5915[123], tmp5915[122], tmp5915[121], tmp5915[120], tmp5915[119], tmp5915[118], tmp5915[117], tmp5915[116], tmp5915[115], tmp5915[114], tmp5915[113], tmp5915[112], tmp5915[111], tmp5915[110], tmp5915[109], tmp5915[108], tmp5915[107], tmp5915[106], tmp5915[105], tmp5915[104], tmp5915[103], tmp5915[102], tmp5915[101], tmp5915[100], tmp5915[99], tmp5915[98], tmp5915[97], tmp5915[96], tmp5915[95], tmp5915[94], tmp5915[93], tmp5915[92], tmp5915[91], tmp5915[90], tmp5915[89], tmp5915[88], tmp5915[87], tmp5915[86], tmp5915[85], tmp5915[84], tmp5915[83], tmp5915[82], tmp5915[81], tmp5915[80], tmp5915[79], tmp5915[78], tmp5915[77], tmp5915[76], tmp5915[75], tmp5915[74], tmp5915[73], tmp5915[72], tmp5915[71], tmp5915[70], tmp5915[69], tmp5915[68], tmp5915[67], tmp5915[66], tmp5915[65], tmp5915[64], tmp5915[63], tmp5915[62], tmp5915[61], tmp5915[60], tmp5915[59], tmp5915[58], tmp5915[57], tmp5915[56], tmp5915[55], tmp5915[54], tmp5915[53], tmp5915[52], tmp5915[51], tmp5915[50], tmp5915[49], tmp5915[48], tmp5915[47], tmp5915[46], tmp5915[45], tmp5915[44], tmp5915[43], tmp5915[42], tmp5915[41], tmp5915[40], tmp5915[39], tmp5915[38], tmp5915[37], tmp5915[36], tmp5915[35], tmp5915[34], tmp5915[33], tmp5915[32], tmp5915[31], tmp5915[30], tmp5915[29], tmp5915[28], tmp5915[27], tmp5915[26], tmp5915[25], tmp5915[24], tmp5915[23], tmp5915[22], tmp5915[21], tmp5915[20], tmp5915[19], tmp5915[18], tmp5915[17], tmp5915[16], tmp5915[15], tmp5915[14], tmp5915[13], tmp5915[12], tmp5915[11], tmp5915[10], tmp5915[9], tmp5915[8], tmp5915[7], tmp5915[6], tmp5915[5], tmp5915[4], tmp5915[3], tmp5915[2], tmp5915[1], tmp5915[0]};
    assign tmp5917 = {tmp5916[255], tmp5916[254], tmp5916[253], tmp5916[252], tmp5916[251], tmp5916[250], tmp5916[249], tmp5916[248], tmp5916[247], tmp5916[246], tmp5916[245], tmp5916[244], tmp5916[243], tmp5916[242], tmp5916[241], tmp5916[240], tmp5916[239], tmp5916[238], tmp5916[237], tmp5916[236], tmp5916[235], tmp5916[234], tmp5916[233], tmp5916[232], tmp5916[231], tmp5916[230], tmp5916[229], tmp5916[228], tmp5916[227], tmp5916[226], tmp5916[225], tmp5916[224], tmp5916[223], tmp5916[222], tmp5916[221], tmp5916[220], tmp5916[219], tmp5916[218], tmp5916[217], tmp5916[216], tmp5916[215], tmp5916[214], tmp5916[213], tmp5916[212], tmp5916[211], tmp5916[210], tmp5916[209], tmp5916[208], tmp5916[207], tmp5916[206], tmp5916[205], tmp5916[204], tmp5916[203], tmp5916[202], tmp5916[201], tmp5916[200], tmp5916[199], tmp5916[198], tmp5916[197], tmp5916[196], tmp5916[195], tmp5916[194], tmp5916[193], tmp5916[192], tmp5916[191], tmp5916[190], tmp5916[189], tmp5916[188], tmp5916[187], tmp5916[186], tmp5916[185], tmp5916[184], tmp5916[183], tmp5916[182], tmp5916[181], tmp5916[180], tmp5916[179], tmp5916[178], tmp5916[177], tmp5916[176], tmp5916[175], tmp5916[174], tmp5916[173], tmp5916[172], tmp5916[171], tmp5916[170], tmp5916[169], tmp5916[168], tmp5916[167], tmp5916[166], tmp5916[165], tmp5916[164], tmp5916[163], tmp5916[162], tmp5916[161], tmp5916[160], tmp5916[159], tmp5916[158], tmp5916[157], tmp5916[156], tmp5916[155], tmp5916[154], tmp5916[153], tmp5916[152], tmp5916[151], tmp5916[150], tmp5916[149], tmp5916[148], tmp5916[147], tmp5916[146], tmp5916[145], tmp5916[144], tmp5916[143], tmp5916[142], tmp5916[141], tmp5916[140], tmp5916[139], tmp5916[138], tmp5916[137], tmp5916[136], tmp5916[135], tmp5916[134], tmp5916[133], tmp5916[132], tmp5916[131], tmp5916[130], tmp5916[129], tmp5916[128], tmp5916[127], tmp5916[126], tmp5916[125], tmp5916[124], tmp5916[123], tmp5916[122], tmp5916[121], tmp5916[120], tmp5916[119], tmp5916[118], tmp5916[117], tmp5916[116], tmp5916[115], tmp5916[114], tmp5916[113], tmp5916[112], tmp5916[111], tmp5916[110], tmp5916[109], tmp5916[108], tmp5916[107], tmp5916[106], tmp5916[105], tmp5916[104], tmp5916[103], tmp5916[102], tmp5916[101], tmp5916[100], tmp5916[99], tmp5916[98], tmp5916[97], tmp5916[96], tmp5916[95], tmp5916[94], tmp5916[93], tmp5916[92], tmp5916[91], tmp5916[90], tmp5916[89], tmp5916[88], tmp5916[87], tmp5916[86], tmp5916[85], tmp5916[84], tmp5916[83], tmp5916[82], tmp5916[81], tmp5916[80], tmp5916[79], tmp5916[78], tmp5916[77], tmp5916[76], tmp5916[75], tmp5916[74], tmp5916[73], tmp5916[72], tmp5916[71], tmp5916[70], tmp5916[69], tmp5916[68], tmp5916[67], tmp5916[66], tmp5916[65], tmp5916[64], tmp5916[63], tmp5916[62], tmp5916[61], tmp5916[60], tmp5916[59], tmp5916[58], tmp5916[57], tmp5916[56], tmp5916[55], tmp5916[54], tmp5916[53], tmp5916[52], tmp5916[51], tmp5916[50], tmp5916[49], tmp5916[48], tmp5916[47], tmp5916[46], tmp5916[45], tmp5916[44], tmp5916[43], tmp5916[42], tmp5916[41], tmp5916[40], tmp5916[39], tmp5916[38], tmp5916[37], tmp5916[36], tmp5916[35], tmp5916[34], tmp5916[33], tmp5916[32], tmp5916[31], tmp5916[30], tmp5916[29], tmp5916[28], tmp5916[27], tmp5916[26], tmp5916[25], tmp5916[24], tmp5916[23], tmp5916[22], tmp5916[21], tmp5916[20], tmp5916[19], tmp5916[18], tmp5916[17], tmp5916[16], tmp5916[15], tmp5916[14], tmp5916[13], tmp5916[12], tmp5916[11], tmp5916[10], tmp5916[9], tmp5916[8], tmp5916[7], tmp5916[6], tmp5916[5], tmp5916[4], tmp5916[3], tmp5916[2], tmp5916[1], tmp5916[0]};
    assign tmp5918 = {const_537_0};
    assign tmp5919 = {tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918, tmp5918};
    assign tmp5920 = {tmp5919, const_537_0};
    assign tmp5921 = {tmp26[255]};
    assign tmp5922 = tmp5920 - tmp26;
    assign tmp5923 = {tmp5922[256]};
    assign tmp5924 = {tmp5920[255]};
    assign tmp5925 = ~tmp5924;
    assign tmp5926 = tmp5923 ^ tmp5925;
    assign tmp5927 = {tmp26[255]};
    assign tmp5928 = ~tmp5927;
    assign tmp5929 = tmp5926 ^ tmp5928;
    assign tmp5930 = {const_538_0};
    assign tmp5931 = {tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930, tmp5930};
    assign tmp5932 = {tmp5931, const_538_0};
    assign tmp5933 = {tmp5908[256]};
    assign tmp5934 = tmp5932 - tmp5908;
    assign tmp5935 = {tmp5934[257]};
    assign tmp5936 = {tmp5932[256]};
    assign tmp5937 = ~tmp5936;
    assign tmp5938 = tmp5935 ^ tmp5937;
    assign tmp5939 = {tmp5908[256]};
    assign tmp5940 = ~tmp5939;
    assign tmp5941 = tmp5938 ^ tmp5940;
    assign tmp5942 = tmp5929 & tmp5941;
    assign tmp5943 = {tmp5917[255]};
    assign tmp5944 = {const_539_0};
    assign tmp5945 = {tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944, tmp5944};
    assign tmp5946 = {tmp5945, const_539_0};
    assign tmp5947 = tmp5917 - tmp5946;
    assign tmp5948 = {tmp5947[256]};
    assign tmp5949 = {tmp5917[255]};
    assign tmp5950 = ~tmp5949;
    assign tmp5951 = tmp5948 ^ tmp5950;
    assign tmp5952 = {tmp5946[255]};
    assign tmp5953 = ~tmp5952;
    assign tmp5954 = tmp5951 ^ tmp5953;
    assign tmp5955 = tmp5917 == tmp5946;
    assign tmp5956 = tmp5954 | tmp5955;
    assign tmp5957 = tmp5942 & tmp5956;
    assign tmp5958 = {tmp26[255]};
    assign tmp5959 = {const_540_0};
    assign tmp5960 = {tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959, tmp5959};
    assign tmp5961 = {tmp5960, const_540_0};
    assign tmp5962 = tmp26 - tmp5961;
    assign tmp5963 = {tmp5962[256]};
    assign tmp5964 = {tmp26[255]};
    assign tmp5965 = ~tmp5964;
    assign tmp5966 = tmp5963 ^ tmp5965;
    assign tmp5967 = {tmp5961[255]};
    assign tmp5968 = ~tmp5967;
    assign tmp5969 = tmp5966 ^ tmp5968;
    assign tmp5970 = {tmp5908[256]};
    assign tmp5971 = {const_541_0};
    assign tmp5972 = {tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971, tmp5971};
    assign tmp5973 = {tmp5972, const_541_0};
    assign tmp5974 = tmp5908 - tmp5973;
    assign tmp5975 = {tmp5974[257]};
    assign tmp5976 = {tmp5908[256]};
    assign tmp5977 = ~tmp5976;
    assign tmp5978 = tmp5975 ^ tmp5977;
    assign tmp5979 = {tmp5973[256]};
    assign tmp5980 = ~tmp5979;
    assign tmp5981 = tmp5978 ^ tmp5980;
    assign tmp5982 = tmp5969 & tmp5981;
    assign tmp5983 = {const_542_0};
    assign tmp5984 = {tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983, tmp5983};
    assign tmp5985 = {tmp5984, const_542_0};
    assign tmp5986 = {tmp5917[255]};
    assign tmp5987 = tmp5985 - tmp5917;
    assign tmp5988 = {tmp5987[256]};
    assign tmp5989 = {tmp5985[255]};
    assign tmp5990 = ~tmp5989;
    assign tmp5991 = tmp5988 ^ tmp5990;
    assign tmp5992 = {tmp5917[255]};
    assign tmp5993 = ~tmp5992;
    assign tmp5994 = tmp5991 ^ tmp5993;
    assign tmp5995 = tmp5985 == tmp5917;
    assign tmp5996 = tmp5994 | tmp5995;
    assign tmp5997 = tmp5982 & tmp5996;
    assign tmp5998 = tmp5957 ? const_543_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp5917;
    assign tmp5999 = tmp5997 ? _ver_out_tmp_49 : tmp5998;
    assign tmp6000 = ~tmp35;
    assign tmp6001 = ~tmp36;
    assign tmp6002 = tmp6000 & tmp6001;
    assign tmp6003 = ~tmp57;
    assign tmp6004 = tmp6002 & tmp6003;
    assign tmp6005 = ~tmp1034;
    assign tmp6006 = tmp6004 & tmp6005;
    assign tmp6007 = tmp6006 & tmp2071;
    assign tmp6008 = ~tmp2583;
    assign tmp6009 = tmp6007 & tmp6008;
    assign tmp6010 = tmp6009 & tmp23;
    assign tmp6011 = ~tmp2627;
    assign tmp6012 = tmp6010 & tmp6011;
    assign tmp6013 = ~tmp2798;
    assign tmp6014 = tmp6012 & tmp6013;
    assign tmp6015 = ~tmp3425;
    assign tmp6016 = tmp6014 & tmp6015;
    assign tmp6017 = ~tmp4020;
    assign tmp6018 = tmp6016 & tmp6017;
    assign tmp6019 = tmp6018 & cfg_speculative_egest;
    assign tmp6020 = ~tmp4511;
    assign tmp6021 = tmp6019 & tmp6020;
    assign tmp6022 = tmp6021 & tmp5688;
    assign tmp6023 = ~tmp35;
    assign tmp6024 = ~tmp36;
    assign tmp6025 = tmp6023 & tmp6024;
    assign tmp6026 = ~tmp57;
    assign tmp6027 = tmp6025 & tmp6026;
    assign tmp6028 = ~tmp1034;
    assign tmp6029 = tmp6027 & tmp6028;
    assign tmp6030 = tmp6029 & tmp2071;
    assign tmp6031 = ~tmp2583;
    assign tmp6032 = tmp6030 & tmp6031;
    assign tmp6033 = tmp6032 & tmp23;
    assign tmp6034 = ~tmp2627;
    assign tmp6035 = tmp6033 & tmp6034;
    assign tmp6036 = ~tmp2798;
    assign tmp6037 = tmp6035 & tmp6036;
    assign tmp6038 = ~tmp3425;
    assign tmp6039 = tmp6037 & tmp6038;
    assign tmp6040 = ~tmp4020;
    assign tmp6041 = tmp6039 & tmp6040;
    assign tmp6042 = tmp6041 & cfg_speculative_egest;
    assign tmp6043 = ~tmp4511;
    assign tmp6044 = tmp6042 & tmp6043;
    assign tmp6045 = tmp6044 & tmp5688;
    assign tmp6046 = _ver_out_tmp_50 == tmp31;
    assign tmp6047 = {const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0, const_547_0};
    assign tmp6048 = {tmp6047, const_546_0};
    assign tmp6049 = tmp6048 - tmp31;
    assign tmp6050 = {const_549_0, const_549_0};
    assign tmp6051 = {tmp6050, const_548_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp6052 = tmp6046 ? tmp6051 : tmp6049;
    assign tmp6053 = {tmp27[255]};
    assign tmp6054 = {tmp6053, tmp6053};
    assign tmp6055 = {tmp6054, tmp27};
    assign tmp6056 = {tmp6052[256]};
    assign tmp6057 = {tmp6056};
    assign tmp6058 = {tmp6057, tmp6052};
    assign tmp6059 = tmp6055 + tmp6058;
    assign tmp6060 = {tmp6059[257], tmp6059[256], tmp6059[255], tmp6059[254], tmp6059[253], tmp6059[252], tmp6059[251], tmp6059[250], tmp6059[249], tmp6059[248], tmp6059[247], tmp6059[246], tmp6059[245], tmp6059[244], tmp6059[243], tmp6059[242], tmp6059[241], tmp6059[240], tmp6059[239], tmp6059[238], tmp6059[237], tmp6059[236], tmp6059[235], tmp6059[234], tmp6059[233], tmp6059[232], tmp6059[231], tmp6059[230], tmp6059[229], tmp6059[228], tmp6059[227], tmp6059[226], tmp6059[225], tmp6059[224], tmp6059[223], tmp6059[222], tmp6059[221], tmp6059[220], tmp6059[219], tmp6059[218], tmp6059[217], tmp6059[216], tmp6059[215], tmp6059[214], tmp6059[213], tmp6059[212], tmp6059[211], tmp6059[210], tmp6059[209], tmp6059[208], tmp6059[207], tmp6059[206], tmp6059[205], tmp6059[204], tmp6059[203], tmp6059[202], tmp6059[201], tmp6059[200], tmp6059[199], tmp6059[198], tmp6059[197], tmp6059[196], tmp6059[195], tmp6059[194], tmp6059[193], tmp6059[192], tmp6059[191], tmp6059[190], tmp6059[189], tmp6059[188], tmp6059[187], tmp6059[186], tmp6059[185], tmp6059[184], tmp6059[183], tmp6059[182], tmp6059[181], tmp6059[180], tmp6059[179], tmp6059[178], tmp6059[177], tmp6059[176], tmp6059[175], tmp6059[174], tmp6059[173], tmp6059[172], tmp6059[171], tmp6059[170], tmp6059[169], tmp6059[168], tmp6059[167], tmp6059[166], tmp6059[165], tmp6059[164], tmp6059[163], tmp6059[162], tmp6059[161], tmp6059[160], tmp6059[159], tmp6059[158], tmp6059[157], tmp6059[156], tmp6059[155], tmp6059[154], tmp6059[153], tmp6059[152], tmp6059[151], tmp6059[150], tmp6059[149], tmp6059[148], tmp6059[147], tmp6059[146], tmp6059[145], tmp6059[144], tmp6059[143], tmp6059[142], tmp6059[141], tmp6059[140], tmp6059[139], tmp6059[138], tmp6059[137], tmp6059[136], tmp6059[135], tmp6059[134], tmp6059[133], tmp6059[132], tmp6059[131], tmp6059[130], tmp6059[129], tmp6059[128], tmp6059[127], tmp6059[126], tmp6059[125], tmp6059[124], tmp6059[123], tmp6059[122], tmp6059[121], tmp6059[120], tmp6059[119], tmp6059[118], tmp6059[117], tmp6059[116], tmp6059[115], tmp6059[114], tmp6059[113], tmp6059[112], tmp6059[111], tmp6059[110], tmp6059[109], tmp6059[108], tmp6059[107], tmp6059[106], tmp6059[105], tmp6059[104], tmp6059[103], tmp6059[102], tmp6059[101], tmp6059[100], tmp6059[99], tmp6059[98], tmp6059[97], tmp6059[96], tmp6059[95], tmp6059[94], tmp6059[93], tmp6059[92], tmp6059[91], tmp6059[90], tmp6059[89], tmp6059[88], tmp6059[87], tmp6059[86], tmp6059[85], tmp6059[84], tmp6059[83], tmp6059[82], tmp6059[81], tmp6059[80], tmp6059[79], tmp6059[78], tmp6059[77], tmp6059[76], tmp6059[75], tmp6059[74], tmp6059[73], tmp6059[72], tmp6059[71], tmp6059[70], tmp6059[69], tmp6059[68], tmp6059[67], tmp6059[66], tmp6059[65], tmp6059[64], tmp6059[63], tmp6059[62], tmp6059[61], tmp6059[60], tmp6059[59], tmp6059[58], tmp6059[57], tmp6059[56], tmp6059[55], tmp6059[54], tmp6059[53], tmp6059[52], tmp6059[51], tmp6059[50], tmp6059[49], tmp6059[48], tmp6059[47], tmp6059[46], tmp6059[45], tmp6059[44], tmp6059[43], tmp6059[42], tmp6059[41], tmp6059[40], tmp6059[39], tmp6059[38], tmp6059[37], tmp6059[36], tmp6059[35], tmp6059[34], tmp6059[33], tmp6059[32], tmp6059[31], tmp6059[30], tmp6059[29], tmp6059[28], tmp6059[27], tmp6059[26], tmp6059[25], tmp6059[24], tmp6059[23], tmp6059[22], tmp6059[21], tmp6059[20], tmp6059[19], tmp6059[18], tmp6059[17], tmp6059[16], tmp6059[15], tmp6059[14], tmp6059[13], tmp6059[12], tmp6059[11], tmp6059[10], tmp6059[9], tmp6059[8], tmp6059[7], tmp6059[6], tmp6059[5], tmp6059[4], tmp6059[3], tmp6059[2], tmp6059[1], tmp6059[0]};
    assign tmp6061 = {tmp6060[255], tmp6060[254], tmp6060[253], tmp6060[252], tmp6060[251], tmp6060[250], tmp6060[249], tmp6060[248], tmp6060[247], tmp6060[246], tmp6060[245], tmp6060[244], tmp6060[243], tmp6060[242], tmp6060[241], tmp6060[240], tmp6060[239], tmp6060[238], tmp6060[237], tmp6060[236], tmp6060[235], tmp6060[234], tmp6060[233], tmp6060[232], tmp6060[231], tmp6060[230], tmp6060[229], tmp6060[228], tmp6060[227], tmp6060[226], tmp6060[225], tmp6060[224], tmp6060[223], tmp6060[222], tmp6060[221], tmp6060[220], tmp6060[219], tmp6060[218], tmp6060[217], tmp6060[216], tmp6060[215], tmp6060[214], tmp6060[213], tmp6060[212], tmp6060[211], tmp6060[210], tmp6060[209], tmp6060[208], tmp6060[207], tmp6060[206], tmp6060[205], tmp6060[204], tmp6060[203], tmp6060[202], tmp6060[201], tmp6060[200], tmp6060[199], tmp6060[198], tmp6060[197], tmp6060[196], tmp6060[195], tmp6060[194], tmp6060[193], tmp6060[192], tmp6060[191], tmp6060[190], tmp6060[189], tmp6060[188], tmp6060[187], tmp6060[186], tmp6060[185], tmp6060[184], tmp6060[183], tmp6060[182], tmp6060[181], tmp6060[180], tmp6060[179], tmp6060[178], tmp6060[177], tmp6060[176], tmp6060[175], tmp6060[174], tmp6060[173], tmp6060[172], tmp6060[171], tmp6060[170], tmp6060[169], tmp6060[168], tmp6060[167], tmp6060[166], tmp6060[165], tmp6060[164], tmp6060[163], tmp6060[162], tmp6060[161], tmp6060[160], tmp6060[159], tmp6060[158], tmp6060[157], tmp6060[156], tmp6060[155], tmp6060[154], tmp6060[153], tmp6060[152], tmp6060[151], tmp6060[150], tmp6060[149], tmp6060[148], tmp6060[147], tmp6060[146], tmp6060[145], tmp6060[144], tmp6060[143], tmp6060[142], tmp6060[141], tmp6060[140], tmp6060[139], tmp6060[138], tmp6060[137], tmp6060[136], tmp6060[135], tmp6060[134], tmp6060[133], tmp6060[132], tmp6060[131], tmp6060[130], tmp6060[129], tmp6060[128], tmp6060[127], tmp6060[126], tmp6060[125], tmp6060[124], tmp6060[123], tmp6060[122], tmp6060[121], tmp6060[120], tmp6060[119], tmp6060[118], tmp6060[117], tmp6060[116], tmp6060[115], tmp6060[114], tmp6060[113], tmp6060[112], tmp6060[111], tmp6060[110], tmp6060[109], tmp6060[108], tmp6060[107], tmp6060[106], tmp6060[105], tmp6060[104], tmp6060[103], tmp6060[102], tmp6060[101], tmp6060[100], tmp6060[99], tmp6060[98], tmp6060[97], tmp6060[96], tmp6060[95], tmp6060[94], tmp6060[93], tmp6060[92], tmp6060[91], tmp6060[90], tmp6060[89], tmp6060[88], tmp6060[87], tmp6060[86], tmp6060[85], tmp6060[84], tmp6060[83], tmp6060[82], tmp6060[81], tmp6060[80], tmp6060[79], tmp6060[78], tmp6060[77], tmp6060[76], tmp6060[75], tmp6060[74], tmp6060[73], tmp6060[72], tmp6060[71], tmp6060[70], tmp6060[69], tmp6060[68], tmp6060[67], tmp6060[66], tmp6060[65], tmp6060[64], tmp6060[63], tmp6060[62], tmp6060[61], tmp6060[60], tmp6060[59], tmp6060[58], tmp6060[57], tmp6060[56], tmp6060[55], tmp6060[54], tmp6060[53], tmp6060[52], tmp6060[51], tmp6060[50], tmp6060[49], tmp6060[48], tmp6060[47], tmp6060[46], tmp6060[45], tmp6060[44], tmp6060[43], tmp6060[42], tmp6060[41], tmp6060[40], tmp6060[39], tmp6060[38], tmp6060[37], tmp6060[36], tmp6060[35], tmp6060[34], tmp6060[33], tmp6060[32], tmp6060[31], tmp6060[30], tmp6060[29], tmp6060[28], tmp6060[27], tmp6060[26], tmp6060[25], tmp6060[24], tmp6060[23], tmp6060[22], tmp6060[21], tmp6060[20], tmp6060[19], tmp6060[18], tmp6060[17], tmp6060[16], tmp6060[15], tmp6060[14], tmp6060[13], tmp6060[12], tmp6060[11], tmp6060[10], tmp6060[9], tmp6060[8], tmp6060[7], tmp6060[6], tmp6060[5], tmp6060[4], tmp6060[3], tmp6060[2], tmp6060[1], tmp6060[0]};
    assign tmp6062 = {const_550_0};
    assign tmp6063 = {tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062, tmp6062};
    assign tmp6064 = {tmp6063, const_550_0};
    assign tmp6065 = {tmp27[255]};
    assign tmp6066 = tmp6064 - tmp27;
    assign tmp6067 = {tmp6066[256]};
    assign tmp6068 = {tmp6064[255]};
    assign tmp6069 = ~tmp6068;
    assign tmp6070 = tmp6067 ^ tmp6069;
    assign tmp6071 = {tmp27[255]};
    assign tmp6072 = ~tmp6071;
    assign tmp6073 = tmp6070 ^ tmp6072;
    assign tmp6074 = {const_551_0};
    assign tmp6075 = {tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074, tmp6074};
    assign tmp6076 = {tmp6075, const_551_0};
    assign tmp6077 = {tmp6052[256]};
    assign tmp6078 = tmp6076 - tmp6052;
    assign tmp6079 = {tmp6078[257]};
    assign tmp6080 = {tmp6076[256]};
    assign tmp6081 = ~tmp6080;
    assign tmp6082 = tmp6079 ^ tmp6081;
    assign tmp6083 = {tmp6052[256]};
    assign tmp6084 = ~tmp6083;
    assign tmp6085 = tmp6082 ^ tmp6084;
    assign tmp6086 = tmp6073 & tmp6085;
    assign tmp6087 = {tmp6061[255]};
    assign tmp6088 = {const_552_0};
    assign tmp6089 = {tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088, tmp6088};
    assign tmp6090 = {tmp6089, const_552_0};
    assign tmp6091 = tmp6061 - tmp6090;
    assign tmp6092 = {tmp6091[256]};
    assign tmp6093 = {tmp6061[255]};
    assign tmp6094 = ~tmp6093;
    assign tmp6095 = tmp6092 ^ tmp6094;
    assign tmp6096 = {tmp6090[255]};
    assign tmp6097 = ~tmp6096;
    assign tmp6098 = tmp6095 ^ tmp6097;
    assign tmp6099 = tmp6061 == tmp6090;
    assign tmp6100 = tmp6098 | tmp6099;
    assign tmp6101 = tmp6086 & tmp6100;
    assign tmp6102 = {tmp27[255]};
    assign tmp6103 = {const_553_0};
    assign tmp6104 = {tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103, tmp6103};
    assign tmp6105 = {tmp6104, const_553_0};
    assign tmp6106 = tmp27 - tmp6105;
    assign tmp6107 = {tmp6106[256]};
    assign tmp6108 = {tmp27[255]};
    assign tmp6109 = ~tmp6108;
    assign tmp6110 = tmp6107 ^ tmp6109;
    assign tmp6111 = {tmp6105[255]};
    assign tmp6112 = ~tmp6111;
    assign tmp6113 = tmp6110 ^ tmp6112;
    assign tmp6114 = {tmp6052[256]};
    assign tmp6115 = {const_554_0};
    assign tmp6116 = {tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115, tmp6115};
    assign tmp6117 = {tmp6116, const_554_0};
    assign tmp6118 = tmp6052 - tmp6117;
    assign tmp6119 = {tmp6118[257]};
    assign tmp6120 = {tmp6052[256]};
    assign tmp6121 = ~tmp6120;
    assign tmp6122 = tmp6119 ^ tmp6121;
    assign tmp6123 = {tmp6117[256]};
    assign tmp6124 = ~tmp6123;
    assign tmp6125 = tmp6122 ^ tmp6124;
    assign tmp6126 = tmp6113 & tmp6125;
    assign tmp6127 = {const_555_0};
    assign tmp6128 = {tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127, tmp6127};
    assign tmp6129 = {tmp6128, const_555_0};
    assign tmp6130 = {tmp6061[255]};
    assign tmp6131 = tmp6129 - tmp6061;
    assign tmp6132 = {tmp6131[256]};
    assign tmp6133 = {tmp6129[255]};
    assign tmp6134 = ~tmp6133;
    assign tmp6135 = tmp6132 ^ tmp6134;
    assign tmp6136 = {tmp6061[255]};
    assign tmp6137 = ~tmp6136;
    assign tmp6138 = tmp6135 ^ tmp6137;
    assign tmp6139 = tmp6129 == tmp6061;
    assign tmp6140 = tmp6138 | tmp6139;
    assign tmp6141 = tmp6126 & tmp6140;
    assign tmp6142 = tmp6101 ? const_556_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp6061;
    assign tmp6143 = tmp6141 ? _ver_out_tmp_56 : tmp6142;
    assign tmp6144 = ~tmp35;
    assign tmp6145 = ~tmp36;
    assign tmp6146 = tmp6144 & tmp6145;
    assign tmp6147 = ~tmp57;
    assign tmp6148 = tmp6146 & tmp6147;
    assign tmp6149 = ~tmp1034;
    assign tmp6150 = tmp6148 & tmp6149;
    assign tmp6151 = tmp6150 & tmp2071;
    assign tmp6152 = ~tmp2583;
    assign tmp6153 = tmp6151 & tmp6152;
    assign tmp6154 = tmp6153 & tmp23;
    assign tmp6155 = ~tmp2627;
    assign tmp6156 = tmp6154 & tmp6155;
    assign tmp6157 = ~tmp2798;
    assign tmp6158 = tmp6156 & tmp6157;
    assign tmp6159 = ~tmp3425;
    assign tmp6160 = tmp6158 & tmp6159;
    assign tmp6161 = ~tmp4020;
    assign tmp6162 = tmp6160 & tmp6161;
    assign tmp6163 = tmp6162 & cfg_speculative_egest;
    assign tmp6164 = ~tmp4511;
    assign tmp6165 = tmp6163 & tmp6164;
    assign tmp6166 = tmp6165 & tmp5688;
    assign tmp6167 = ~tmp35;
    assign tmp6168 = ~tmp36;
    assign tmp6169 = tmp6167 & tmp6168;
    assign tmp6170 = ~tmp57;
    assign tmp6171 = tmp6169 & tmp6170;
    assign tmp6172 = ~tmp1034;
    assign tmp6173 = tmp6171 & tmp6172;
    assign tmp6174 = tmp6173 & tmp2071;
    assign tmp6175 = ~tmp2583;
    assign tmp6176 = tmp6174 & tmp6175;
    assign tmp6177 = tmp6176 & tmp23;
    assign tmp6178 = ~tmp2627;
    assign tmp6179 = tmp6177 & tmp6178;
    assign tmp6180 = ~tmp2798;
    assign tmp6181 = tmp6179 & tmp6180;
    assign tmp6182 = ~tmp3425;
    assign tmp6183 = tmp6181 & tmp6182;
    assign tmp6184 = ~tmp4020;
    assign tmp6185 = tmp6183 & tmp6184;
    assign tmp6186 = tmp6185 & cfg_speculative_egest;
    assign tmp6187 = ~tmp4511;
    assign tmp6188 = tmp6186 & tmp6187;
    assign tmp6189 = tmp6188 & tmp5688;
    assign tmp6190 = _ver_out_tmp_57 == tmp32;
    assign tmp6191 = {const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0, const_560_0};
    assign tmp6192 = {tmp6191, const_559_0};
    assign tmp6193 = tmp6192 - tmp32;
    assign tmp6194 = {const_562_0, const_562_0};
    assign tmp6195 = {tmp6194, const_561_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp6196 = tmp6190 ? tmp6195 : tmp6193;
    assign tmp6197 = {tmp28[255]};
    assign tmp6198 = {tmp6197, tmp6197};
    assign tmp6199 = {tmp6198, tmp28};
    assign tmp6200 = {tmp6196[256]};
    assign tmp6201 = {tmp6200};
    assign tmp6202 = {tmp6201, tmp6196};
    assign tmp6203 = tmp6199 + tmp6202;
    assign tmp6204 = {tmp6203[257], tmp6203[256], tmp6203[255], tmp6203[254], tmp6203[253], tmp6203[252], tmp6203[251], tmp6203[250], tmp6203[249], tmp6203[248], tmp6203[247], tmp6203[246], tmp6203[245], tmp6203[244], tmp6203[243], tmp6203[242], tmp6203[241], tmp6203[240], tmp6203[239], tmp6203[238], tmp6203[237], tmp6203[236], tmp6203[235], tmp6203[234], tmp6203[233], tmp6203[232], tmp6203[231], tmp6203[230], tmp6203[229], tmp6203[228], tmp6203[227], tmp6203[226], tmp6203[225], tmp6203[224], tmp6203[223], tmp6203[222], tmp6203[221], tmp6203[220], tmp6203[219], tmp6203[218], tmp6203[217], tmp6203[216], tmp6203[215], tmp6203[214], tmp6203[213], tmp6203[212], tmp6203[211], tmp6203[210], tmp6203[209], tmp6203[208], tmp6203[207], tmp6203[206], tmp6203[205], tmp6203[204], tmp6203[203], tmp6203[202], tmp6203[201], tmp6203[200], tmp6203[199], tmp6203[198], tmp6203[197], tmp6203[196], tmp6203[195], tmp6203[194], tmp6203[193], tmp6203[192], tmp6203[191], tmp6203[190], tmp6203[189], tmp6203[188], tmp6203[187], tmp6203[186], tmp6203[185], tmp6203[184], tmp6203[183], tmp6203[182], tmp6203[181], tmp6203[180], tmp6203[179], tmp6203[178], tmp6203[177], tmp6203[176], tmp6203[175], tmp6203[174], tmp6203[173], tmp6203[172], tmp6203[171], tmp6203[170], tmp6203[169], tmp6203[168], tmp6203[167], tmp6203[166], tmp6203[165], tmp6203[164], tmp6203[163], tmp6203[162], tmp6203[161], tmp6203[160], tmp6203[159], tmp6203[158], tmp6203[157], tmp6203[156], tmp6203[155], tmp6203[154], tmp6203[153], tmp6203[152], tmp6203[151], tmp6203[150], tmp6203[149], tmp6203[148], tmp6203[147], tmp6203[146], tmp6203[145], tmp6203[144], tmp6203[143], tmp6203[142], tmp6203[141], tmp6203[140], tmp6203[139], tmp6203[138], tmp6203[137], tmp6203[136], tmp6203[135], tmp6203[134], tmp6203[133], tmp6203[132], tmp6203[131], tmp6203[130], tmp6203[129], tmp6203[128], tmp6203[127], tmp6203[126], tmp6203[125], tmp6203[124], tmp6203[123], tmp6203[122], tmp6203[121], tmp6203[120], tmp6203[119], tmp6203[118], tmp6203[117], tmp6203[116], tmp6203[115], tmp6203[114], tmp6203[113], tmp6203[112], tmp6203[111], tmp6203[110], tmp6203[109], tmp6203[108], tmp6203[107], tmp6203[106], tmp6203[105], tmp6203[104], tmp6203[103], tmp6203[102], tmp6203[101], tmp6203[100], tmp6203[99], tmp6203[98], tmp6203[97], tmp6203[96], tmp6203[95], tmp6203[94], tmp6203[93], tmp6203[92], tmp6203[91], tmp6203[90], tmp6203[89], tmp6203[88], tmp6203[87], tmp6203[86], tmp6203[85], tmp6203[84], tmp6203[83], tmp6203[82], tmp6203[81], tmp6203[80], tmp6203[79], tmp6203[78], tmp6203[77], tmp6203[76], tmp6203[75], tmp6203[74], tmp6203[73], tmp6203[72], tmp6203[71], tmp6203[70], tmp6203[69], tmp6203[68], tmp6203[67], tmp6203[66], tmp6203[65], tmp6203[64], tmp6203[63], tmp6203[62], tmp6203[61], tmp6203[60], tmp6203[59], tmp6203[58], tmp6203[57], tmp6203[56], tmp6203[55], tmp6203[54], tmp6203[53], tmp6203[52], tmp6203[51], tmp6203[50], tmp6203[49], tmp6203[48], tmp6203[47], tmp6203[46], tmp6203[45], tmp6203[44], tmp6203[43], tmp6203[42], tmp6203[41], tmp6203[40], tmp6203[39], tmp6203[38], tmp6203[37], tmp6203[36], tmp6203[35], tmp6203[34], tmp6203[33], tmp6203[32], tmp6203[31], tmp6203[30], tmp6203[29], tmp6203[28], tmp6203[27], tmp6203[26], tmp6203[25], tmp6203[24], tmp6203[23], tmp6203[22], tmp6203[21], tmp6203[20], tmp6203[19], tmp6203[18], tmp6203[17], tmp6203[16], tmp6203[15], tmp6203[14], tmp6203[13], tmp6203[12], tmp6203[11], tmp6203[10], tmp6203[9], tmp6203[8], tmp6203[7], tmp6203[6], tmp6203[5], tmp6203[4], tmp6203[3], tmp6203[2], tmp6203[1], tmp6203[0]};
    assign tmp6205 = {tmp6204[255], tmp6204[254], tmp6204[253], tmp6204[252], tmp6204[251], tmp6204[250], tmp6204[249], tmp6204[248], tmp6204[247], tmp6204[246], tmp6204[245], tmp6204[244], tmp6204[243], tmp6204[242], tmp6204[241], tmp6204[240], tmp6204[239], tmp6204[238], tmp6204[237], tmp6204[236], tmp6204[235], tmp6204[234], tmp6204[233], tmp6204[232], tmp6204[231], tmp6204[230], tmp6204[229], tmp6204[228], tmp6204[227], tmp6204[226], tmp6204[225], tmp6204[224], tmp6204[223], tmp6204[222], tmp6204[221], tmp6204[220], tmp6204[219], tmp6204[218], tmp6204[217], tmp6204[216], tmp6204[215], tmp6204[214], tmp6204[213], tmp6204[212], tmp6204[211], tmp6204[210], tmp6204[209], tmp6204[208], tmp6204[207], tmp6204[206], tmp6204[205], tmp6204[204], tmp6204[203], tmp6204[202], tmp6204[201], tmp6204[200], tmp6204[199], tmp6204[198], tmp6204[197], tmp6204[196], tmp6204[195], tmp6204[194], tmp6204[193], tmp6204[192], tmp6204[191], tmp6204[190], tmp6204[189], tmp6204[188], tmp6204[187], tmp6204[186], tmp6204[185], tmp6204[184], tmp6204[183], tmp6204[182], tmp6204[181], tmp6204[180], tmp6204[179], tmp6204[178], tmp6204[177], tmp6204[176], tmp6204[175], tmp6204[174], tmp6204[173], tmp6204[172], tmp6204[171], tmp6204[170], tmp6204[169], tmp6204[168], tmp6204[167], tmp6204[166], tmp6204[165], tmp6204[164], tmp6204[163], tmp6204[162], tmp6204[161], tmp6204[160], tmp6204[159], tmp6204[158], tmp6204[157], tmp6204[156], tmp6204[155], tmp6204[154], tmp6204[153], tmp6204[152], tmp6204[151], tmp6204[150], tmp6204[149], tmp6204[148], tmp6204[147], tmp6204[146], tmp6204[145], tmp6204[144], tmp6204[143], tmp6204[142], tmp6204[141], tmp6204[140], tmp6204[139], tmp6204[138], tmp6204[137], tmp6204[136], tmp6204[135], tmp6204[134], tmp6204[133], tmp6204[132], tmp6204[131], tmp6204[130], tmp6204[129], tmp6204[128], tmp6204[127], tmp6204[126], tmp6204[125], tmp6204[124], tmp6204[123], tmp6204[122], tmp6204[121], tmp6204[120], tmp6204[119], tmp6204[118], tmp6204[117], tmp6204[116], tmp6204[115], tmp6204[114], tmp6204[113], tmp6204[112], tmp6204[111], tmp6204[110], tmp6204[109], tmp6204[108], tmp6204[107], tmp6204[106], tmp6204[105], tmp6204[104], tmp6204[103], tmp6204[102], tmp6204[101], tmp6204[100], tmp6204[99], tmp6204[98], tmp6204[97], tmp6204[96], tmp6204[95], tmp6204[94], tmp6204[93], tmp6204[92], tmp6204[91], tmp6204[90], tmp6204[89], tmp6204[88], tmp6204[87], tmp6204[86], tmp6204[85], tmp6204[84], tmp6204[83], tmp6204[82], tmp6204[81], tmp6204[80], tmp6204[79], tmp6204[78], tmp6204[77], tmp6204[76], tmp6204[75], tmp6204[74], tmp6204[73], tmp6204[72], tmp6204[71], tmp6204[70], tmp6204[69], tmp6204[68], tmp6204[67], tmp6204[66], tmp6204[65], tmp6204[64], tmp6204[63], tmp6204[62], tmp6204[61], tmp6204[60], tmp6204[59], tmp6204[58], tmp6204[57], tmp6204[56], tmp6204[55], tmp6204[54], tmp6204[53], tmp6204[52], tmp6204[51], tmp6204[50], tmp6204[49], tmp6204[48], tmp6204[47], tmp6204[46], tmp6204[45], tmp6204[44], tmp6204[43], tmp6204[42], tmp6204[41], tmp6204[40], tmp6204[39], tmp6204[38], tmp6204[37], tmp6204[36], tmp6204[35], tmp6204[34], tmp6204[33], tmp6204[32], tmp6204[31], tmp6204[30], tmp6204[29], tmp6204[28], tmp6204[27], tmp6204[26], tmp6204[25], tmp6204[24], tmp6204[23], tmp6204[22], tmp6204[21], tmp6204[20], tmp6204[19], tmp6204[18], tmp6204[17], tmp6204[16], tmp6204[15], tmp6204[14], tmp6204[13], tmp6204[12], tmp6204[11], tmp6204[10], tmp6204[9], tmp6204[8], tmp6204[7], tmp6204[6], tmp6204[5], tmp6204[4], tmp6204[3], tmp6204[2], tmp6204[1], tmp6204[0]};
    assign tmp6206 = {const_563_0};
    assign tmp6207 = {tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206, tmp6206};
    assign tmp6208 = {tmp6207, const_563_0};
    assign tmp6209 = {tmp28[255]};
    assign tmp6210 = tmp6208 - tmp28;
    assign tmp6211 = {tmp6210[256]};
    assign tmp6212 = {tmp6208[255]};
    assign tmp6213 = ~tmp6212;
    assign tmp6214 = tmp6211 ^ tmp6213;
    assign tmp6215 = {tmp28[255]};
    assign tmp6216 = ~tmp6215;
    assign tmp6217 = tmp6214 ^ tmp6216;
    assign tmp6218 = {const_564_0};
    assign tmp6219 = {tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218, tmp6218};
    assign tmp6220 = {tmp6219, const_564_0};
    assign tmp6221 = {tmp6196[256]};
    assign tmp6222 = tmp6220 - tmp6196;
    assign tmp6223 = {tmp6222[257]};
    assign tmp6224 = {tmp6220[256]};
    assign tmp6225 = ~tmp6224;
    assign tmp6226 = tmp6223 ^ tmp6225;
    assign tmp6227 = {tmp6196[256]};
    assign tmp6228 = ~tmp6227;
    assign tmp6229 = tmp6226 ^ tmp6228;
    assign tmp6230 = tmp6217 & tmp6229;
    assign tmp6231 = {tmp6205[255]};
    assign tmp6232 = {const_565_0};
    assign tmp6233 = {tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232, tmp6232};
    assign tmp6234 = {tmp6233, const_565_0};
    assign tmp6235 = tmp6205 - tmp6234;
    assign tmp6236 = {tmp6235[256]};
    assign tmp6237 = {tmp6205[255]};
    assign tmp6238 = ~tmp6237;
    assign tmp6239 = tmp6236 ^ tmp6238;
    assign tmp6240 = {tmp6234[255]};
    assign tmp6241 = ~tmp6240;
    assign tmp6242 = tmp6239 ^ tmp6241;
    assign tmp6243 = tmp6205 == tmp6234;
    assign tmp6244 = tmp6242 | tmp6243;
    assign tmp6245 = tmp6230 & tmp6244;
    assign tmp6246 = {tmp28[255]};
    assign tmp6247 = {const_566_0};
    assign tmp6248 = {tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247, tmp6247};
    assign tmp6249 = {tmp6248, const_566_0};
    assign tmp6250 = tmp28 - tmp6249;
    assign tmp6251 = {tmp6250[256]};
    assign tmp6252 = {tmp28[255]};
    assign tmp6253 = ~tmp6252;
    assign tmp6254 = tmp6251 ^ tmp6253;
    assign tmp6255 = {tmp6249[255]};
    assign tmp6256 = ~tmp6255;
    assign tmp6257 = tmp6254 ^ tmp6256;
    assign tmp6258 = {tmp6196[256]};
    assign tmp6259 = {const_567_0};
    assign tmp6260 = {tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259, tmp6259};
    assign tmp6261 = {tmp6260, const_567_0};
    assign tmp6262 = tmp6196 - tmp6261;
    assign tmp6263 = {tmp6262[257]};
    assign tmp6264 = {tmp6196[256]};
    assign tmp6265 = ~tmp6264;
    assign tmp6266 = tmp6263 ^ tmp6265;
    assign tmp6267 = {tmp6261[256]};
    assign tmp6268 = ~tmp6267;
    assign tmp6269 = tmp6266 ^ tmp6268;
    assign tmp6270 = tmp6257 & tmp6269;
    assign tmp6271 = {const_568_0};
    assign tmp6272 = {tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271, tmp6271};
    assign tmp6273 = {tmp6272, const_568_0};
    assign tmp6274 = {tmp6205[255]};
    assign tmp6275 = tmp6273 - tmp6205;
    assign tmp6276 = {tmp6275[256]};
    assign tmp6277 = {tmp6273[255]};
    assign tmp6278 = ~tmp6277;
    assign tmp6279 = tmp6276 ^ tmp6278;
    assign tmp6280 = {tmp6205[255]};
    assign tmp6281 = ~tmp6280;
    assign tmp6282 = tmp6279 ^ tmp6281;
    assign tmp6283 = tmp6273 == tmp6205;
    assign tmp6284 = tmp6282 | tmp6283;
    assign tmp6285 = tmp6270 & tmp6284;
    assign tmp6286 = tmp6245 ? const_569_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp6205;
    assign tmp6287 = tmp6285 ? _ver_out_tmp_3 : tmp6286;
    assign tmp6288 = ~tmp35;
    assign tmp6289 = ~tmp36;
    assign tmp6290 = tmp6288 & tmp6289;
    assign tmp6291 = ~tmp57;
    assign tmp6292 = tmp6290 & tmp6291;
    assign tmp6293 = ~tmp1034;
    assign tmp6294 = tmp6292 & tmp6293;
    assign tmp6295 = tmp6294 & tmp2071;
    assign tmp6296 = ~tmp2583;
    assign tmp6297 = tmp6295 & tmp6296;
    assign tmp6298 = tmp6297 & tmp23;
    assign tmp6299 = ~tmp2627;
    assign tmp6300 = tmp6298 & tmp6299;
    assign tmp6301 = ~tmp2798;
    assign tmp6302 = tmp6300 & tmp6301;
    assign tmp6303 = ~tmp3425;
    assign tmp6304 = tmp6302 & tmp6303;
    assign tmp6305 = ~tmp4020;
    assign tmp6306 = tmp6304 & tmp6305;
    assign tmp6307 = tmp6306 & cfg_speculative_egest;
    assign tmp6308 = ~tmp4511;
    assign tmp6309 = tmp6307 & tmp6308;
    assign tmp6310 = tmp6309 & tmp5688;
    assign tmp6311 = ~tmp35;
    assign tmp6312 = ~tmp36;
    assign tmp6313 = tmp6311 & tmp6312;
    assign tmp6314 = ~tmp57;
    assign tmp6315 = tmp6313 & tmp6314;
    assign tmp6316 = ~tmp1034;
    assign tmp6317 = tmp6315 & tmp6316;
    assign tmp6318 = tmp6317 & tmp2071;
    assign tmp6319 = ~tmp2583;
    assign tmp6320 = tmp6318 & tmp6319;
    assign tmp6321 = tmp6320 & tmp23;
    assign tmp6322 = ~tmp2627;
    assign tmp6323 = tmp6321 & tmp6322;
    assign tmp6324 = ~tmp2798;
    assign tmp6325 = tmp6323 & tmp6324;
    assign tmp6326 = ~tmp3425;
    assign tmp6327 = tmp6325 & tmp6326;
    assign tmp6328 = ~tmp4020;
    assign tmp6329 = tmp6327 & tmp6328;
    assign tmp6330 = tmp6329 & cfg_speculative_egest;
    assign tmp6331 = ~tmp4511;
    assign tmp6332 = tmp6330 & tmp6331;
    assign tmp6333 = ~tmp5688;
    assign tmp6334 = tmp6332 & tmp6333;
    assign tmp6335 = ~tmp35;
    assign tmp6336 = ~tmp36;
    assign tmp6337 = tmp6335 & tmp6336;
    assign tmp6338 = ~tmp57;
    assign tmp6339 = tmp6337 & tmp6338;
    assign tmp6340 = ~tmp1034;
    assign tmp6341 = tmp6339 & tmp6340;
    assign tmp6342 = tmp6341 & tmp2071;
    assign tmp6343 = ~tmp2583;
    assign tmp6344 = tmp6342 & tmp6343;
    assign tmp6345 = tmp6344 & tmp23;
    assign tmp6346 = ~tmp2627;
    assign tmp6347 = tmp6345 & tmp6346;
    assign tmp6348 = ~tmp2798;
    assign tmp6349 = tmp6347 & tmp6348;
    assign tmp6350 = ~tmp3425;
    assign tmp6351 = tmp6349 & tmp6350;
    assign tmp6352 = ~tmp4020;
    assign tmp6353 = tmp6351 & tmp6352;
    assign tmp6354 = tmp6353 & cfg_speculative_egest;
    assign tmp6355 = ~tmp4511;
    assign tmp6356 = tmp6354 & tmp6355;
    assign tmp6357 = ~tmp5688;
    assign tmp6358 = tmp6356 & tmp6357;
    assign tmp6359 = ~tmp35;
    assign tmp6360 = ~tmp36;
    assign tmp6361 = tmp6359 & tmp6360;
    assign tmp6362 = ~tmp57;
    assign tmp6363 = tmp6361 & tmp6362;
    assign tmp6364 = ~tmp1034;
    assign tmp6365 = tmp6363 & tmp6364;
    assign tmp6366 = tmp6365 & tmp2071;
    assign tmp6367 = ~tmp2583;
    assign tmp6368 = tmp6366 & tmp6367;
    assign tmp6369 = tmp6368 & tmp23;
    assign tmp6370 = ~tmp2627;
    assign tmp6371 = tmp6369 & tmp6370;
    assign tmp6372 = ~tmp2798;
    assign tmp6373 = tmp6371 & tmp6372;
    assign tmp6374 = ~tmp3425;
    assign tmp6375 = tmp6373 & tmp6374;
    assign tmp6376 = ~tmp4020;
    assign tmp6377 = tmp6375 & tmp6376;
    assign tmp6378 = ~cfg_speculative_egest;
    assign tmp6379 = tmp6377 & tmp6378;
    assign tmp6380 = ~tmp35;
    assign tmp6381 = ~tmp36;
    assign tmp6382 = tmp6380 & tmp6381;
    assign tmp6383 = ~tmp57;
    assign tmp6384 = tmp6382 & tmp6383;
    assign tmp6385 = ~tmp1034;
    assign tmp6386 = tmp6384 & tmp6385;
    assign tmp6387 = tmp6386 & tmp2071;
    assign tmp6388 = ~tmp2583;
    assign tmp6389 = tmp6387 & tmp6388;
    assign tmp6390 = tmp6389 & tmp23;
    assign tmp6391 = ~tmp2627;
    assign tmp6392 = tmp6390 & tmp6391;
    assign tmp6393 = ~tmp2798;
    assign tmp6394 = tmp6392 & tmp6393;
    assign tmp6395 = ~tmp3425;
    assign tmp6396 = tmp6394 & tmp6395;
    assign tmp6397 = ~tmp4020;
    assign tmp6398 = tmp6396 & tmp6397;
    assign tmp6399 = ~cfg_speculative_egest;
    assign tmp6400 = tmp6398 & tmp6399;
    assign tmp6401 = {tmp11[255]};
    assign tmp6402 = {const_575_0};
    assign tmp6403 = {tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402, tmp6402};
    assign tmp6404 = {tmp6403, const_575_0};
    assign tmp6405 = tmp11 - tmp6404;
    assign tmp6406 = {tmp6405[256]};
    assign tmp6407 = {tmp11[255]};
    assign tmp6408 = ~tmp6407;
    assign tmp6409 = tmp6406 ^ tmp6408;
    assign tmp6410 = {tmp6404[255]};
    assign tmp6411 = ~tmp6410;
    assign tmp6412 = tmp6409 ^ tmp6411;
    assign tmp6413 = tmp11 == _ver_out_tmp_5;
    assign tmp6414 = {const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0, const_578_0};
    assign tmp6415 = {tmp6414, const_577_0};
    assign tmp6416 = tmp6415 - tmp11;
    assign tmp6417 = {const_580_0, const_580_0};
    assign tmp6418 = {tmp6417, const_579_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp6419 = tmp6413 ? tmp6418 : tmp6416;
    assign tmp6420 = {const_581_0};
    assign tmp6421 = {tmp6420, tmp11};
    assign tmp6422 = tmp6412 ? tmp6421 : tmp6419;
    assign tmp6423 = {tmp15[255]};
    assign tmp6424 = {const_582_0};
    assign tmp6425 = {tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424, tmp6424};
    assign tmp6426 = {tmp6425, const_582_0};
    assign tmp6427 = tmp15 - tmp6426;
    assign tmp6428 = {tmp6427[256]};
    assign tmp6429 = {tmp15[255]};
    assign tmp6430 = ~tmp6429;
    assign tmp6431 = tmp6428 ^ tmp6430;
    assign tmp6432 = {tmp6426[255]};
    assign tmp6433 = ~tmp6432;
    assign tmp6434 = tmp6431 ^ tmp6433;
    assign tmp6435 = tmp15 == _ver_out_tmp_6;
    assign tmp6436 = {const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0, const_585_0};
    assign tmp6437 = {tmp6436, const_584_0};
    assign tmp6438 = tmp6437 - tmp15;
    assign tmp6439 = {const_587_0, const_587_0};
    assign tmp6440 = {tmp6439, const_586_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp6441 = tmp6435 ? tmp6440 : tmp6438;
    assign tmp6442 = {const_588_0};
    assign tmp6443 = {tmp6442, tmp15};
    assign tmp6444 = tmp6434 ? tmp6443 : tmp6441;
    assign tmp6445 = {tmp6422[256]};
    assign tmp6446 = {tmp6444[256]};
    assign tmp6447 = tmp6422 - tmp6444;
    assign tmp6448 = {tmp6447[257]};
    assign tmp6449 = {tmp6422[256]};
    assign tmp6450 = ~tmp6449;
    assign tmp6451 = tmp6448 ^ tmp6450;
    assign tmp6452 = {tmp6444[256]};
    assign tmp6453 = ~tmp6452;
    assign tmp6454 = tmp6451 ^ tmp6453;
    assign tmp6455 = {tmp12[255]};
    assign tmp6456 = {const_589_0};
    assign tmp6457 = {tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456, tmp6456};
    assign tmp6458 = {tmp6457, const_589_0};
    assign tmp6459 = tmp12 - tmp6458;
    assign tmp6460 = {tmp6459[256]};
    assign tmp6461 = {tmp12[255]};
    assign tmp6462 = ~tmp6461;
    assign tmp6463 = tmp6460 ^ tmp6462;
    assign tmp6464 = {tmp6458[255]};
    assign tmp6465 = ~tmp6464;
    assign tmp6466 = tmp6463 ^ tmp6465;
    assign tmp6467 = tmp12 == _ver_out_tmp_8;
    assign tmp6468 = {const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0, const_592_0};
    assign tmp6469 = {tmp6468, const_591_0};
    assign tmp6470 = tmp6469 - tmp12;
    assign tmp6471 = {const_594_0, const_594_0};
    assign tmp6472 = {tmp6471, const_593_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp6473 = tmp6467 ? tmp6472 : tmp6470;
    assign tmp6474 = {const_595_0};
    assign tmp6475 = {tmp6474, tmp12};
    assign tmp6476 = tmp6466 ? tmp6475 : tmp6473;
    assign tmp6477 = {tmp16[255]};
    assign tmp6478 = {const_596_0};
    assign tmp6479 = {tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478, tmp6478};
    assign tmp6480 = {tmp6479, const_596_0};
    assign tmp6481 = tmp16 - tmp6480;
    assign tmp6482 = {tmp6481[256]};
    assign tmp6483 = {tmp16[255]};
    assign tmp6484 = ~tmp6483;
    assign tmp6485 = tmp6482 ^ tmp6484;
    assign tmp6486 = {tmp6480[255]};
    assign tmp6487 = ~tmp6486;
    assign tmp6488 = tmp6485 ^ tmp6487;
    assign tmp6489 = tmp16 == _ver_out_tmp_51;
    assign tmp6490 = {const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0, const_599_0};
    assign tmp6491 = {tmp6490, const_598_0};
    assign tmp6492 = tmp6491 - tmp16;
    assign tmp6493 = {const_601_0, const_601_0};
    assign tmp6494 = {tmp6493, const_600_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp6495 = tmp6489 ? tmp6494 : tmp6492;
    assign tmp6496 = {const_602_0};
    assign tmp6497 = {tmp6496, tmp16};
    assign tmp6498 = tmp6488 ? tmp6497 : tmp6495;
    assign tmp6499 = {tmp6476[256]};
    assign tmp6500 = {tmp6498[256]};
    assign tmp6501 = tmp6476 - tmp6498;
    assign tmp6502 = {tmp6501[257]};
    assign tmp6503 = {tmp6476[256]};
    assign tmp6504 = ~tmp6503;
    assign tmp6505 = tmp6502 ^ tmp6504;
    assign tmp6506 = {tmp6498[256]};
    assign tmp6507 = ~tmp6506;
    assign tmp6508 = tmp6505 ^ tmp6507;
    assign tmp6509 = tmp6454 & tmp6508;
    assign tmp6510 = {tmp13[255]};
    assign tmp6511 = {const_603_0};
    assign tmp6512 = {tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511, tmp6511};
    assign tmp6513 = {tmp6512, const_603_0};
    assign tmp6514 = tmp13 - tmp6513;
    assign tmp6515 = {tmp6514[256]};
    assign tmp6516 = {tmp13[255]};
    assign tmp6517 = ~tmp6516;
    assign tmp6518 = tmp6515 ^ tmp6517;
    assign tmp6519 = {tmp6513[255]};
    assign tmp6520 = ~tmp6519;
    assign tmp6521 = tmp6518 ^ tmp6520;
    assign tmp6522 = tmp13 == _ver_out_tmp_11;
    assign tmp6523 = {const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0, const_606_0};
    assign tmp6524 = {tmp6523, const_605_0};
    assign tmp6525 = tmp6524 - tmp13;
    assign tmp6526 = {const_608_0, const_608_0};
    assign tmp6527 = {tmp6526, const_607_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp6528 = tmp6522 ? tmp6527 : tmp6525;
    assign tmp6529 = {const_609_0};
    assign tmp6530 = {tmp6529, tmp13};
    assign tmp6531 = tmp6521 ? tmp6530 : tmp6528;
    assign tmp6532 = {tmp17[255]};
    assign tmp6533 = {const_610_0};
    assign tmp6534 = {tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533, tmp6533};
    assign tmp6535 = {tmp6534, const_610_0};
    assign tmp6536 = tmp17 - tmp6535;
    assign tmp6537 = {tmp6536[256]};
    assign tmp6538 = {tmp17[255]};
    assign tmp6539 = ~tmp6538;
    assign tmp6540 = tmp6537 ^ tmp6539;
    assign tmp6541 = {tmp6535[255]};
    assign tmp6542 = ~tmp6541;
    assign tmp6543 = tmp6540 ^ tmp6542;
    assign tmp6544 = tmp17 == _ver_out_tmp_13;
    assign tmp6545 = {const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0, const_613_0};
    assign tmp6546 = {tmp6545, const_612_0};
    assign tmp6547 = tmp6546 - tmp17;
    assign tmp6548 = {const_615_0, const_615_0};
    assign tmp6549 = {tmp6548, const_614_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp6550 = tmp6544 ? tmp6549 : tmp6547;
    assign tmp6551 = {const_616_0};
    assign tmp6552 = {tmp6551, tmp17};
    assign tmp6553 = tmp6543 ? tmp6552 : tmp6550;
    assign tmp6554 = {tmp6531[256]};
    assign tmp6555 = {tmp6553[256]};
    assign tmp6556 = tmp6531 - tmp6553;
    assign tmp6557 = {tmp6556[257]};
    assign tmp6558 = {tmp6531[256]};
    assign tmp6559 = ~tmp6558;
    assign tmp6560 = tmp6557 ^ tmp6559;
    assign tmp6561 = {tmp6553[256]};
    assign tmp6562 = ~tmp6561;
    assign tmp6563 = tmp6560 ^ tmp6562;
    assign tmp6564 = tmp6509 & tmp6563;
    assign tmp6565 = {tmp14[255]};
    assign tmp6566 = {const_617_0};
    assign tmp6567 = {tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566, tmp6566};
    assign tmp6568 = {tmp6567, const_617_0};
    assign tmp6569 = tmp14 - tmp6568;
    assign tmp6570 = {tmp6569[256]};
    assign tmp6571 = {tmp14[255]};
    assign tmp6572 = ~tmp6571;
    assign tmp6573 = tmp6570 ^ tmp6572;
    assign tmp6574 = {tmp6568[255]};
    assign tmp6575 = ~tmp6574;
    assign tmp6576 = tmp6573 ^ tmp6575;
    assign tmp6577 = tmp14 == _ver_out_tmp_17;
    assign tmp6578 = {const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0, const_620_0};
    assign tmp6579 = {tmp6578, const_619_0};
    assign tmp6580 = tmp6579 - tmp14;
    assign tmp6581 = {const_622_0, const_622_0};
    assign tmp6582 = {tmp6581, const_621_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp6583 = tmp6577 ? tmp6582 : tmp6580;
    assign tmp6584 = {const_623_0};
    assign tmp6585 = {tmp6584, tmp14};
    assign tmp6586 = tmp6576 ? tmp6585 : tmp6583;
    assign tmp6587 = {tmp18[255]};
    assign tmp6588 = {const_624_0};
    assign tmp6589 = {tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588, tmp6588};
    assign tmp6590 = {tmp6589, const_624_0};
    assign tmp6591 = tmp18 - tmp6590;
    assign tmp6592 = {tmp6591[256]};
    assign tmp6593 = {tmp18[255]};
    assign tmp6594 = ~tmp6593;
    assign tmp6595 = tmp6592 ^ tmp6594;
    assign tmp6596 = {tmp6590[255]};
    assign tmp6597 = ~tmp6596;
    assign tmp6598 = tmp6595 ^ tmp6597;
    assign tmp6599 = tmp18 == _ver_out_tmp_20;
    assign tmp6600 = {const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0, const_627_0};
    assign tmp6601 = {tmp6600, const_626_0};
    assign tmp6602 = tmp6601 - tmp18;
    assign tmp6603 = {const_629_0, const_629_0};
    assign tmp6604 = {tmp6603, const_628_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp6605 = tmp6599 ? tmp6604 : tmp6602;
    assign tmp6606 = {const_630_0};
    assign tmp6607 = {tmp6606, tmp18};
    assign tmp6608 = tmp6598 ? tmp6607 : tmp6605;
    assign tmp6609 = {tmp6586[256]};
    assign tmp6610 = {tmp6608[256]};
    assign tmp6611 = tmp6586 - tmp6608;
    assign tmp6612 = {tmp6611[257]};
    assign tmp6613 = {tmp6586[256]};
    assign tmp6614 = ~tmp6613;
    assign tmp6615 = tmp6612 ^ tmp6614;
    assign tmp6616 = {tmp6608[256]};
    assign tmp6617 = ~tmp6616;
    assign tmp6618 = tmp6615 ^ tmp6617;
    assign tmp6619 = tmp6564 & tmp6618;
    assign tmp6620 = ~tmp35;
    assign tmp6621 = ~tmp36;
    assign tmp6622 = tmp6620 & tmp6621;
    assign tmp6623 = ~tmp57;
    assign tmp6624 = tmp6622 & tmp6623;
    assign tmp6625 = ~tmp1034;
    assign tmp6626 = tmp6624 & tmp6625;
    assign tmp6627 = tmp6626 & tmp2071;
    assign tmp6628 = ~tmp2583;
    assign tmp6629 = tmp6627 & tmp6628;
    assign tmp6630 = ~tmp23;
    assign tmp6631 = tmp6629 & tmp6630;
    assign tmp6632 = tmp6631 & cfg_speculative_egest;
    assign tmp6633 = tmp6632 & tmp6619;
    assign tmp6634 = ~tmp35;
    assign tmp6635 = ~tmp36;
    assign tmp6636 = tmp6634 & tmp6635;
    assign tmp6637 = ~tmp57;
    assign tmp6638 = tmp6636 & tmp6637;
    assign tmp6639 = ~tmp1034;
    assign tmp6640 = tmp6638 & tmp6639;
    assign tmp6641 = tmp6640 & tmp2071;
    assign tmp6642 = ~tmp2583;
    assign tmp6643 = tmp6641 & tmp6642;
    assign tmp6644 = ~tmp23;
    assign tmp6645 = tmp6643 & tmp6644;
    assign tmp6646 = tmp6645 & cfg_speculative_egest;
    assign tmp6647 = tmp6646 & tmp6619;
    assign tmp6648 = ~tmp35;
    assign tmp6649 = ~tmp36;
    assign tmp6650 = tmp6648 & tmp6649;
    assign tmp6651 = ~tmp57;
    assign tmp6652 = tmp6650 & tmp6651;
    assign tmp6653 = ~tmp1034;
    assign tmp6654 = tmp6652 & tmp6653;
    assign tmp6655 = tmp6654 & tmp2071;
    assign tmp6656 = ~tmp2583;
    assign tmp6657 = tmp6655 & tmp6656;
    assign tmp6658 = ~tmp23;
    assign tmp6659 = tmp6657 & tmp6658;
    assign tmp6660 = tmp6659 & cfg_speculative_egest;
    assign tmp6661 = tmp6660 & tmp6619;
    assign tmp6662 = ~tmp35;
    assign tmp6663 = ~tmp36;
    assign tmp6664 = tmp6662 & tmp6663;
    assign tmp6665 = ~tmp57;
    assign tmp6666 = tmp6664 & tmp6665;
    assign tmp6667 = ~tmp1034;
    assign tmp6668 = tmp6666 & tmp6667;
    assign tmp6669 = tmp6668 & tmp2071;
    assign tmp6670 = ~tmp2583;
    assign tmp6671 = tmp6669 & tmp6670;
    assign tmp6672 = ~tmp23;
    assign tmp6673 = tmp6671 & tmp6672;
    assign tmp6674 = tmp6673 & cfg_speculative_egest;
    assign tmp6675 = tmp6674 & tmp6619;
    assign tmp6676 = ~tmp35;
    assign tmp6677 = ~tmp36;
    assign tmp6678 = tmp6676 & tmp6677;
    assign tmp6679 = ~tmp57;
    assign tmp6680 = tmp6678 & tmp6679;
    assign tmp6681 = ~tmp1034;
    assign tmp6682 = tmp6680 & tmp6681;
    assign tmp6683 = tmp6682 & tmp2071;
    assign tmp6684 = ~tmp2583;
    assign tmp6685 = tmp6683 & tmp6684;
    assign tmp6686 = ~tmp23;
    assign tmp6687 = tmp6685 & tmp6686;
    assign tmp6688 = tmp6687 & cfg_speculative_egest;
    assign tmp6689 = tmp6688 & tmp6619;
    assign tmp6690 = ~tmp35;
    assign tmp6691 = ~tmp36;
    assign tmp6692 = tmp6690 & tmp6691;
    assign tmp6693 = ~tmp57;
    assign tmp6694 = tmp6692 & tmp6693;
    assign tmp6695 = ~tmp1034;
    assign tmp6696 = tmp6694 & tmp6695;
    assign tmp6697 = tmp6696 & tmp2071;
    assign tmp6698 = ~tmp2583;
    assign tmp6699 = tmp6697 & tmp6698;
    assign tmp6700 = ~tmp23;
    assign tmp6701 = tmp6699 & tmp6700;
    assign tmp6702 = tmp6701 & cfg_speculative_egest;
    assign tmp6703 = tmp6702 & tmp6619;
    assign tmp6704 = ~tmp35;
    assign tmp6705 = ~tmp36;
    assign tmp6706 = tmp6704 & tmp6705;
    assign tmp6707 = ~tmp57;
    assign tmp6708 = tmp6706 & tmp6707;
    assign tmp6709 = ~tmp1034;
    assign tmp6710 = tmp6708 & tmp6709;
    assign tmp6711 = tmp6710 & tmp2071;
    assign tmp6712 = ~tmp2583;
    assign tmp6713 = tmp6711 & tmp6712;
    assign tmp6714 = ~tmp23;
    assign tmp6715 = tmp6713 & tmp6714;
    assign tmp6716 = tmp6715 & cfg_speculative_egest;
    assign tmp6717 = tmp6716 & tmp6619;
    assign tmp6718 = ~tmp35;
    assign tmp6719 = ~tmp36;
    assign tmp6720 = tmp6718 & tmp6719;
    assign tmp6721 = ~tmp57;
    assign tmp6722 = tmp6720 & tmp6721;
    assign tmp6723 = ~tmp1034;
    assign tmp6724 = tmp6722 & tmp6723;
    assign tmp6725 = tmp6724 & tmp2071;
    assign tmp6726 = ~tmp2583;
    assign tmp6727 = tmp6725 & tmp6726;
    assign tmp6728 = ~tmp23;
    assign tmp6729 = tmp6727 & tmp6728;
    assign tmp6730 = tmp6729 & cfg_speculative_egest;
    assign tmp6731 = tmp6730 & tmp6619;
    assign tmp6732 = ~tmp35;
    assign tmp6733 = ~tmp36;
    assign tmp6734 = tmp6732 & tmp6733;
    assign tmp6735 = ~tmp57;
    assign tmp6736 = tmp6734 & tmp6735;
    assign tmp6737 = ~tmp1034;
    assign tmp6738 = tmp6736 & tmp6737;
    assign tmp6739 = tmp6738 & tmp2071;
    assign tmp6740 = ~tmp2583;
    assign tmp6741 = tmp6739 & tmp6740;
    assign tmp6742 = ~tmp23;
    assign tmp6743 = tmp6741 & tmp6742;
    assign tmp6744 = tmp6743 & cfg_speculative_egest;
    assign tmp6745 = tmp6744 & tmp6619;
    assign tmp6746 = ~tmp35;
    assign tmp6747 = ~tmp36;
    assign tmp6748 = tmp6746 & tmp6747;
    assign tmp6749 = ~tmp57;
    assign tmp6750 = tmp6748 & tmp6749;
    assign tmp6751 = ~tmp1034;
    assign tmp6752 = tmp6750 & tmp6751;
    assign tmp6753 = tmp6752 & tmp2071;
    assign tmp6754 = ~tmp2583;
    assign tmp6755 = tmp6753 & tmp6754;
    assign tmp6756 = ~tmp23;
    assign tmp6757 = tmp6755 & tmp6756;
    assign tmp6758 = tmp6757 & cfg_speculative_egest;
    assign tmp6759 = tmp6758 & tmp6619;
    assign tmp6760 = {tmp11[255]};
    assign tmp6761 = {const_633_0};
    assign tmp6762 = {tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761, tmp6761};
    assign tmp6763 = {tmp6762, const_633_0};
    assign tmp6764 = tmp11 - tmp6763;
    assign tmp6765 = {tmp6764[256]};
    assign tmp6766 = {tmp11[255]};
    assign tmp6767 = ~tmp6766;
    assign tmp6768 = tmp6765 ^ tmp6767;
    assign tmp6769 = {tmp6763[255]};
    assign tmp6770 = ~tmp6769;
    assign tmp6771 = tmp6768 ^ tmp6770;
    assign tmp6772 = tmp11 == _ver_out_tmp_25;
    assign tmp6773 = {const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0, const_636_0};
    assign tmp6774 = {tmp6773, const_635_0};
    assign tmp6775 = tmp6774 - tmp11;
    assign tmp6776 = {const_638_0, const_638_0};
    assign tmp6777 = {tmp6776, const_637_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp6778 = tmp6772 ? tmp6777 : tmp6775;
    assign tmp6779 = {const_639_0};
    assign tmp6780 = {tmp6779, tmp11};
    assign tmp6781 = tmp6771 ? tmp6780 : tmp6778;
    assign tmp6782 = {tmp6781[256], tmp6781[255], tmp6781[254], tmp6781[253], tmp6781[252], tmp6781[251], tmp6781[250], tmp6781[249], tmp6781[248], tmp6781[247], tmp6781[246], tmp6781[245], tmp6781[244], tmp6781[243], tmp6781[242], tmp6781[241], tmp6781[240], tmp6781[239], tmp6781[238], tmp6781[237], tmp6781[236], tmp6781[235], tmp6781[234], tmp6781[233], tmp6781[232], tmp6781[231], tmp6781[230], tmp6781[229], tmp6781[228], tmp6781[227], tmp6781[226], tmp6781[225], tmp6781[224], tmp6781[223], tmp6781[222], tmp6781[221], tmp6781[220], tmp6781[219], tmp6781[218], tmp6781[217], tmp6781[216], tmp6781[215], tmp6781[214], tmp6781[213], tmp6781[212], tmp6781[211], tmp6781[210], tmp6781[209], tmp6781[208], tmp6781[207], tmp6781[206], tmp6781[205], tmp6781[204], tmp6781[203], tmp6781[202], tmp6781[201], tmp6781[200], tmp6781[199], tmp6781[198], tmp6781[197], tmp6781[196], tmp6781[195], tmp6781[194], tmp6781[193], tmp6781[192], tmp6781[191], tmp6781[190], tmp6781[189], tmp6781[188], tmp6781[187], tmp6781[186], tmp6781[185], tmp6781[184], tmp6781[183], tmp6781[182], tmp6781[181], tmp6781[180], tmp6781[179], tmp6781[178], tmp6781[177], tmp6781[176], tmp6781[175], tmp6781[174], tmp6781[173], tmp6781[172], tmp6781[171], tmp6781[170], tmp6781[169], tmp6781[168], tmp6781[167], tmp6781[166], tmp6781[165], tmp6781[164], tmp6781[163], tmp6781[162], tmp6781[161], tmp6781[160], tmp6781[159], tmp6781[158], tmp6781[157], tmp6781[156], tmp6781[155], tmp6781[154], tmp6781[153], tmp6781[152], tmp6781[151], tmp6781[150], tmp6781[149], tmp6781[148], tmp6781[147], tmp6781[146], tmp6781[145], tmp6781[144], tmp6781[143], tmp6781[142], tmp6781[141], tmp6781[140], tmp6781[139], tmp6781[138], tmp6781[137], tmp6781[136], tmp6781[135], tmp6781[134], tmp6781[133], tmp6781[132], tmp6781[131], tmp6781[130], tmp6781[129], tmp6781[128], tmp6781[127], tmp6781[126], tmp6781[125], tmp6781[124], tmp6781[123], tmp6781[122], tmp6781[121], tmp6781[120], tmp6781[119], tmp6781[118], tmp6781[117], tmp6781[116], tmp6781[115], tmp6781[114], tmp6781[113], tmp6781[112], tmp6781[111], tmp6781[110], tmp6781[109], tmp6781[108], tmp6781[107], tmp6781[106], tmp6781[105], tmp6781[104], tmp6781[103], tmp6781[102], tmp6781[101], tmp6781[100], tmp6781[99], tmp6781[98], tmp6781[97], tmp6781[96], tmp6781[95], tmp6781[94], tmp6781[93], tmp6781[92], tmp6781[91], tmp6781[90], tmp6781[89], tmp6781[88], tmp6781[87], tmp6781[86], tmp6781[85], tmp6781[84], tmp6781[83], tmp6781[82], tmp6781[81], tmp6781[80], tmp6781[79], tmp6781[78], tmp6781[77], tmp6781[76], tmp6781[75], tmp6781[74], tmp6781[73], tmp6781[72], tmp6781[71], tmp6781[70], tmp6781[69], tmp6781[68], tmp6781[67], tmp6781[66], tmp6781[65], tmp6781[64], tmp6781[63], tmp6781[62], tmp6781[61], tmp6781[60], tmp6781[59], tmp6781[58], tmp6781[57], tmp6781[56], tmp6781[55], tmp6781[54], tmp6781[53], tmp6781[52], tmp6781[51], tmp6781[50], tmp6781[49], tmp6781[48], tmp6781[47], tmp6781[46], tmp6781[45], tmp6781[44], tmp6781[43], tmp6781[42], tmp6781[41], tmp6781[40], tmp6781[39], tmp6781[38], tmp6781[37], tmp6781[36], tmp6781[35], tmp6781[34], tmp6781[33], tmp6781[32], tmp6781[31], tmp6781[30], tmp6781[29], tmp6781[28], tmp6781[27], tmp6781[26], tmp6781[25], tmp6781[24], tmp6781[23], tmp6781[22], tmp6781[21], tmp6781[20], tmp6781[19], tmp6781[18], tmp6781[17], tmp6781[16], tmp6781[15], tmp6781[14], tmp6781[13], tmp6781[12], tmp6781[11], tmp6781[10], tmp6781[9], tmp6781[8], tmp6781[7], tmp6781[6], tmp6781[5], tmp6781[4], tmp6781[3], tmp6781[2], tmp6781[1]};
    assign tmp6783 = {tmp6782[255]};
    assign tmp6784 = {tmp6783};
    assign tmp6785 = {tmp6784, tmp6782};
    assign tmp6786 = {tmp15[255]};
    assign tmp6787 = {const_640_0};
    assign tmp6788 = {tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787, tmp6787};
    assign tmp6789 = {tmp6788, const_640_0};
    assign tmp6790 = tmp15 - tmp6789;
    assign tmp6791 = {tmp6790[256]};
    assign tmp6792 = {tmp15[255]};
    assign tmp6793 = ~tmp6792;
    assign tmp6794 = tmp6791 ^ tmp6793;
    assign tmp6795 = {tmp6789[255]};
    assign tmp6796 = ~tmp6795;
    assign tmp6797 = tmp6794 ^ tmp6796;
    assign tmp6798 = tmp15 == _ver_out_tmp_27;
    assign tmp6799 = {const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0, const_643_0};
    assign tmp6800 = {tmp6799, const_642_0};
    assign tmp6801 = tmp6800 - tmp15;
    assign tmp6802 = {const_645_0, const_645_0};
    assign tmp6803 = {tmp6802, const_644_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp6804 = tmp6798 ? tmp6803 : tmp6801;
    assign tmp6805 = {const_646_0};
    assign tmp6806 = {tmp6805, tmp15};
    assign tmp6807 = tmp6797 ? tmp6806 : tmp6804;
    assign tmp6808 = {tmp6785[256]};
    assign tmp6809 = {tmp6807[256]};
    assign tmp6810 = tmp6807 - tmp6785;
    assign tmp6811 = {tmp6810[257]};
    assign tmp6812 = {tmp6785[256]};
    assign tmp6813 = ~tmp6812;
    assign tmp6814 = tmp6811 ^ tmp6813;
    assign tmp6815 = {tmp6807[256]};
    assign tmp6816 = ~tmp6815;
    assign tmp6817 = tmp6814 ^ tmp6816;
    assign tmp6818 = tmp6785 == tmp6807;
    assign tmp6819 = tmp6817 | tmp6818;
    assign tmp6820 = tmp19 & tmp6819;
    assign tmp6821 = {tmp12[255]};
    assign tmp6822 = {const_647_0};
    assign tmp6823 = {tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822, tmp6822};
    assign tmp6824 = {tmp6823, const_647_0};
    assign tmp6825 = tmp12 - tmp6824;
    assign tmp6826 = {tmp6825[256]};
    assign tmp6827 = {tmp12[255]};
    assign tmp6828 = ~tmp6827;
    assign tmp6829 = tmp6826 ^ tmp6828;
    assign tmp6830 = {tmp6824[255]};
    assign tmp6831 = ~tmp6830;
    assign tmp6832 = tmp6829 ^ tmp6831;
    assign tmp6833 = tmp12 == _ver_out_tmp_29;
    assign tmp6834 = {const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0, const_650_0};
    assign tmp6835 = {tmp6834, const_649_0};
    assign tmp6836 = tmp6835 - tmp12;
    assign tmp6837 = {const_652_0, const_652_0};
    assign tmp6838 = {tmp6837, const_651_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp6839 = tmp6833 ? tmp6838 : tmp6836;
    assign tmp6840 = {const_653_0};
    assign tmp6841 = {tmp6840, tmp12};
    assign tmp6842 = tmp6832 ? tmp6841 : tmp6839;
    assign tmp6843 = {tmp6842[256], tmp6842[255], tmp6842[254], tmp6842[253], tmp6842[252], tmp6842[251], tmp6842[250], tmp6842[249], tmp6842[248], tmp6842[247], tmp6842[246], tmp6842[245], tmp6842[244], tmp6842[243], tmp6842[242], tmp6842[241], tmp6842[240], tmp6842[239], tmp6842[238], tmp6842[237], tmp6842[236], tmp6842[235], tmp6842[234], tmp6842[233], tmp6842[232], tmp6842[231], tmp6842[230], tmp6842[229], tmp6842[228], tmp6842[227], tmp6842[226], tmp6842[225], tmp6842[224], tmp6842[223], tmp6842[222], tmp6842[221], tmp6842[220], tmp6842[219], tmp6842[218], tmp6842[217], tmp6842[216], tmp6842[215], tmp6842[214], tmp6842[213], tmp6842[212], tmp6842[211], tmp6842[210], tmp6842[209], tmp6842[208], tmp6842[207], tmp6842[206], tmp6842[205], tmp6842[204], tmp6842[203], tmp6842[202], tmp6842[201], tmp6842[200], tmp6842[199], tmp6842[198], tmp6842[197], tmp6842[196], tmp6842[195], tmp6842[194], tmp6842[193], tmp6842[192], tmp6842[191], tmp6842[190], tmp6842[189], tmp6842[188], tmp6842[187], tmp6842[186], tmp6842[185], tmp6842[184], tmp6842[183], tmp6842[182], tmp6842[181], tmp6842[180], tmp6842[179], tmp6842[178], tmp6842[177], tmp6842[176], tmp6842[175], tmp6842[174], tmp6842[173], tmp6842[172], tmp6842[171], tmp6842[170], tmp6842[169], tmp6842[168], tmp6842[167], tmp6842[166], tmp6842[165], tmp6842[164], tmp6842[163], tmp6842[162], tmp6842[161], tmp6842[160], tmp6842[159], tmp6842[158], tmp6842[157], tmp6842[156], tmp6842[155], tmp6842[154], tmp6842[153], tmp6842[152], tmp6842[151], tmp6842[150], tmp6842[149], tmp6842[148], tmp6842[147], tmp6842[146], tmp6842[145], tmp6842[144], tmp6842[143], tmp6842[142], tmp6842[141], tmp6842[140], tmp6842[139], tmp6842[138], tmp6842[137], tmp6842[136], tmp6842[135], tmp6842[134], tmp6842[133], tmp6842[132], tmp6842[131], tmp6842[130], tmp6842[129], tmp6842[128], tmp6842[127], tmp6842[126], tmp6842[125], tmp6842[124], tmp6842[123], tmp6842[122], tmp6842[121], tmp6842[120], tmp6842[119], tmp6842[118], tmp6842[117], tmp6842[116], tmp6842[115], tmp6842[114], tmp6842[113], tmp6842[112], tmp6842[111], tmp6842[110], tmp6842[109], tmp6842[108], tmp6842[107], tmp6842[106], tmp6842[105], tmp6842[104], tmp6842[103], tmp6842[102], tmp6842[101], tmp6842[100], tmp6842[99], tmp6842[98], tmp6842[97], tmp6842[96], tmp6842[95], tmp6842[94], tmp6842[93], tmp6842[92], tmp6842[91], tmp6842[90], tmp6842[89], tmp6842[88], tmp6842[87], tmp6842[86], tmp6842[85], tmp6842[84], tmp6842[83], tmp6842[82], tmp6842[81], tmp6842[80], tmp6842[79], tmp6842[78], tmp6842[77], tmp6842[76], tmp6842[75], tmp6842[74], tmp6842[73], tmp6842[72], tmp6842[71], tmp6842[70], tmp6842[69], tmp6842[68], tmp6842[67], tmp6842[66], tmp6842[65], tmp6842[64], tmp6842[63], tmp6842[62], tmp6842[61], tmp6842[60], tmp6842[59], tmp6842[58], tmp6842[57], tmp6842[56], tmp6842[55], tmp6842[54], tmp6842[53], tmp6842[52], tmp6842[51], tmp6842[50], tmp6842[49], tmp6842[48], tmp6842[47], tmp6842[46], tmp6842[45], tmp6842[44], tmp6842[43], tmp6842[42], tmp6842[41], tmp6842[40], tmp6842[39], tmp6842[38], tmp6842[37], tmp6842[36], tmp6842[35], tmp6842[34], tmp6842[33], tmp6842[32], tmp6842[31], tmp6842[30], tmp6842[29], tmp6842[28], tmp6842[27], tmp6842[26], tmp6842[25], tmp6842[24], tmp6842[23], tmp6842[22], tmp6842[21], tmp6842[20], tmp6842[19], tmp6842[18], tmp6842[17], tmp6842[16], tmp6842[15], tmp6842[14], tmp6842[13], tmp6842[12], tmp6842[11], tmp6842[10], tmp6842[9], tmp6842[8], tmp6842[7], tmp6842[6], tmp6842[5], tmp6842[4], tmp6842[3], tmp6842[2], tmp6842[1]};
    assign tmp6844 = {tmp6843[255]};
    assign tmp6845 = {tmp6844};
    assign tmp6846 = {tmp6845, tmp6843};
    assign tmp6847 = {tmp16[255]};
    assign tmp6848 = {const_654_0};
    assign tmp6849 = {tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848, tmp6848};
    assign tmp6850 = {tmp6849, const_654_0};
    assign tmp6851 = tmp16 - tmp6850;
    assign tmp6852 = {tmp6851[256]};
    assign tmp6853 = {tmp16[255]};
    assign tmp6854 = ~tmp6853;
    assign tmp6855 = tmp6852 ^ tmp6854;
    assign tmp6856 = {tmp6850[255]};
    assign tmp6857 = ~tmp6856;
    assign tmp6858 = tmp6855 ^ tmp6857;
    assign tmp6859 = tmp16 == _ver_out_tmp_32;
    assign tmp6860 = {const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0, const_657_0};
    assign tmp6861 = {tmp6860, const_656_0};
    assign tmp6862 = tmp6861 - tmp16;
    assign tmp6863 = {const_659_0, const_659_0};
    assign tmp6864 = {tmp6863, const_658_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp6865 = tmp6859 ? tmp6864 : tmp6862;
    assign tmp6866 = {const_660_0};
    assign tmp6867 = {tmp6866, tmp16};
    assign tmp6868 = tmp6858 ? tmp6867 : tmp6865;
    assign tmp6869 = {tmp6846[256]};
    assign tmp6870 = {tmp6868[256]};
    assign tmp6871 = tmp6868 - tmp6846;
    assign tmp6872 = {tmp6871[257]};
    assign tmp6873 = {tmp6846[256]};
    assign tmp6874 = ~tmp6873;
    assign tmp6875 = tmp6872 ^ tmp6874;
    assign tmp6876 = {tmp6868[256]};
    assign tmp6877 = ~tmp6876;
    assign tmp6878 = tmp6875 ^ tmp6877;
    assign tmp6879 = tmp6846 == tmp6868;
    assign tmp6880 = tmp6878 | tmp6879;
    assign tmp6881 = tmp6820 & tmp6880;
    assign tmp6882 = {tmp13[255]};
    assign tmp6883 = {const_661_0};
    assign tmp6884 = {tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883, tmp6883};
    assign tmp6885 = {tmp6884, const_661_0};
    assign tmp6886 = tmp13 - tmp6885;
    assign tmp6887 = {tmp6886[256]};
    assign tmp6888 = {tmp13[255]};
    assign tmp6889 = ~tmp6888;
    assign tmp6890 = tmp6887 ^ tmp6889;
    assign tmp6891 = {tmp6885[255]};
    assign tmp6892 = ~tmp6891;
    assign tmp6893 = tmp6890 ^ tmp6892;
    assign tmp6894 = tmp13 == _ver_out_tmp_36;
    assign tmp6895 = {const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0, const_664_0};
    assign tmp6896 = {tmp6895, const_663_0};
    assign tmp6897 = tmp6896 - tmp13;
    assign tmp6898 = {const_666_0, const_666_0};
    assign tmp6899 = {tmp6898, const_665_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp6900 = tmp6894 ? tmp6899 : tmp6897;
    assign tmp6901 = {const_667_0};
    assign tmp6902 = {tmp6901, tmp13};
    assign tmp6903 = tmp6893 ? tmp6902 : tmp6900;
    assign tmp6904 = {tmp6903[256], tmp6903[255], tmp6903[254], tmp6903[253], tmp6903[252], tmp6903[251], tmp6903[250], tmp6903[249], tmp6903[248], tmp6903[247], tmp6903[246], tmp6903[245], tmp6903[244], tmp6903[243], tmp6903[242], tmp6903[241], tmp6903[240], tmp6903[239], tmp6903[238], tmp6903[237], tmp6903[236], tmp6903[235], tmp6903[234], tmp6903[233], tmp6903[232], tmp6903[231], tmp6903[230], tmp6903[229], tmp6903[228], tmp6903[227], tmp6903[226], tmp6903[225], tmp6903[224], tmp6903[223], tmp6903[222], tmp6903[221], tmp6903[220], tmp6903[219], tmp6903[218], tmp6903[217], tmp6903[216], tmp6903[215], tmp6903[214], tmp6903[213], tmp6903[212], tmp6903[211], tmp6903[210], tmp6903[209], tmp6903[208], tmp6903[207], tmp6903[206], tmp6903[205], tmp6903[204], tmp6903[203], tmp6903[202], tmp6903[201], tmp6903[200], tmp6903[199], tmp6903[198], tmp6903[197], tmp6903[196], tmp6903[195], tmp6903[194], tmp6903[193], tmp6903[192], tmp6903[191], tmp6903[190], tmp6903[189], tmp6903[188], tmp6903[187], tmp6903[186], tmp6903[185], tmp6903[184], tmp6903[183], tmp6903[182], tmp6903[181], tmp6903[180], tmp6903[179], tmp6903[178], tmp6903[177], tmp6903[176], tmp6903[175], tmp6903[174], tmp6903[173], tmp6903[172], tmp6903[171], tmp6903[170], tmp6903[169], tmp6903[168], tmp6903[167], tmp6903[166], tmp6903[165], tmp6903[164], tmp6903[163], tmp6903[162], tmp6903[161], tmp6903[160], tmp6903[159], tmp6903[158], tmp6903[157], tmp6903[156], tmp6903[155], tmp6903[154], tmp6903[153], tmp6903[152], tmp6903[151], tmp6903[150], tmp6903[149], tmp6903[148], tmp6903[147], tmp6903[146], tmp6903[145], tmp6903[144], tmp6903[143], tmp6903[142], tmp6903[141], tmp6903[140], tmp6903[139], tmp6903[138], tmp6903[137], tmp6903[136], tmp6903[135], tmp6903[134], tmp6903[133], tmp6903[132], tmp6903[131], tmp6903[130], tmp6903[129], tmp6903[128], tmp6903[127], tmp6903[126], tmp6903[125], tmp6903[124], tmp6903[123], tmp6903[122], tmp6903[121], tmp6903[120], tmp6903[119], tmp6903[118], tmp6903[117], tmp6903[116], tmp6903[115], tmp6903[114], tmp6903[113], tmp6903[112], tmp6903[111], tmp6903[110], tmp6903[109], tmp6903[108], tmp6903[107], tmp6903[106], tmp6903[105], tmp6903[104], tmp6903[103], tmp6903[102], tmp6903[101], tmp6903[100], tmp6903[99], tmp6903[98], tmp6903[97], tmp6903[96], tmp6903[95], tmp6903[94], tmp6903[93], tmp6903[92], tmp6903[91], tmp6903[90], tmp6903[89], tmp6903[88], tmp6903[87], tmp6903[86], tmp6903[85], tmp6903[84], tmp6903[83], tmp6903[82], tmp6903[81], tmp6903[80], tmp6903[79], tmp6903[78], tmp6903[77], tmp6903[76], tmp6903[75], tmp6903[74], tmp6903[73], tmp6903[72], tmp6903[71], tmp6903[70], tmp6903[69], tmp6903[68], tmp6903[67], tmp6903[66], tmp6903[65], tmp6903[64], tmp6903[63], tmp6903[62], tmp6903[61], tmp6903[60], tmp6903[59], tmp6903[58], tmp6903[57], tmp6903[56], tmp6903[55], tmp6903[54], tmp6903[53], tmp6903[52], tmp6903[51], tmp6903[50], tmp6903[49], tmp6903[48], tmp6903[47], tmp6903[46], tmp6903[45], tmp6903[44], tmp6903[43], tmp6903[42], tmp6903[41], tmp6903[40], tmp6903[39], tmp6903[38], tmp6903[37], tmp6903[36], tmp6903[35], tmp6903[34], tmp6903[33], tmp6903[32], tmp6903[31], tmp6903[30], tmp6903[29], tmp6903[28], tmp6903[27], tmp6903[26], tmp6903[25], tmp6903[24], tmp6903[23], tmp6903[22], tmp6903[21], tmp6903[20], tmp6903[19], tmp6903[18], tmp6903[17], tmp6903[16], tmp6903[15], tmp6903[14], tmp6903[13], tmp6903[12], tmp6903[11], tmp6903[10], tmp6903[9], tmp6903[8], tmp6903[7], tmp6903[6], tmp6903[5], tmp6903[4], tmp6903[3], tmp6903[2], tmp6903[1]};
    assign tmp6905 = {tmp6904[255]};
    assign tmp6906 = {tmp6905};
    assign tmp6907 = {tmp6906, tmp6904};
    assign tmp6908 = {tmp17[255]};
    assign tmp6909 = {const_668_0};
    assign tmp6910 = {tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909, tmp6909};
    assign tmp6911 = {tmp6910, const_668_0};
    assign tmp6912 = tmp17 - tmp6911;
    assign tmp6913 = {tmp6912[256]};
    assign tmp6914 = {tmp17[255]};
    assign tmp6915 = ~tmp6914;
    assign tmp6916 = tmp6913 ^ tmp6915;
    assign tmp6917 = {tmp6911[255]};
    assign tmp6918 = ~tmp6917;
    assign tmp6919 = tmp6916 ^ tmp6918;
    assign tmp6920 = tmp17 == _ver_out_tmp_68;
    assign tmp6921 = {const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0, const_671_0};
    assign tmp6922 = {tmp6921, const_670_0};
    assign tmp6923 = tmp6922 - tmp17;
    assign tmp6924 = {const_673_0, const_673_0};
    assign tmp6925 = {tmp6924, const_672_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp6926 = tmp6920 ? tmp6925 : tmp6923;
    assign tmp6927 = {const_674_0};
    assign tmp6928 = {tmp6927, tmp17};
    assign tmp6929 = tmp6919 ? tmp6928 : tmp6926;
    assign tmp6930 = {tmp6907[256]};
    assign tmp6931 = {tmp6929[256]};
    assign tmp6932 = tmp6929 - tmp6907;
    assign tmp6933 = {tmp6932[257]};
    assign tmp6934 = {tmp6907[256]};
    assign tmp6935 = ~tmp6934;
    assign tmp6936 = tmp6933 ^ tmp6935;
    assign tmp6937 = {tmp6929[256]};
    assign tmp6938 = ~tmp6937;
    assign tmp6939 = tmp6936 ^ tmp6938;
    assign tmp6940 = tmp6907 == tmp6929;
    assign tmp6941 = tmp6939 | tmp6940;
    assign tmp6942 = tmp6881 & tmp6941;
    assign tmp6943 = {tmp14[255]};
    assign tmp6944 = {const_675_0};
    assign tmp6945 = {tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944, tmp6944};
    assign tmp6946 = {tmp6945, const_675_0};
    assign tmp6947 = tmp14 - tmp6946;
    assign tmp6948 = {tmp6947[256]};
    assign tmp6949 = {tmp14[255]};
    assign tmp6950 = ~tmp6949;
    assign tmp6951 = tmp6948 ^ tmp6950;
    assign tmp6952 = {tmp6946[255]};
    assign tmp6953 = ~tmp6952;
    assign tmp6954 = tmp6951 ^ tmp6953;
    assign tmp6955 = tmp14 == _ver_out_tmp_43;
    assign tmp6956 = {const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0, const_678_0};
    assign tmp6957 = {tmp6956, const_677_0};
    assign tmp6958 = tmp6957 - tmp14;
    assign tmp6959 = {const_680_0, const_680_0};
    assign tmp6960 = {tmp6959, const_679_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp6961 = tmp6955 ? tmp6960 : tmp6958;
    assign tmp6962 = {const_681_0};
    assign tmp6963 = {tmp6962, tmp14};
    assign tmp6964 = tmp6954 ? tmp6963 : tmp6961;
    assign tmp6965 = {tmp6964[256], tmp6964[255], tmp6964[254], tmp6964[253], tmp6964[252], tmp6964[251], tmp6964[250], tmp6964[249], tmp6964[248], tmp6964[247], tmp6964[246], tmp6964[245], tmp6964[244], tmp6964[243], tmp6964[242], tmp6964[241], tmp6964[240], tmp6964[239], tmp6964[238], tmp6964[237], tmp6964[236], tmp6964[235], tmp6964[234], tmp6964[233], tmp6964[232], tmp6964[231], tmp6964[230], tmp6964[229], tmp6964[228], tmp6964[227], tmp6964[226], tmp6964[225], tmp6964[224], tmp6964[223], tmp6964[222], tmp6964[221], tmp6964[220], tmp6964[219], tmp6964[218], tmp6964[217], tmp6964[216], tmp6964[215], tmp6964[214], tmp6964[213], tmp6964[212], tmp6964[211], tmp6964[210], tmp6964[209], tmp6964[208], tmp6964[207], tmp6964[206], tmp6964[205], tmp6964[204], tmp6964[203], tmp6964[202], tmp6964[201], tmp6964[200], tmp6964[199], tmp6964[198], tmp6964[197], tmp6964[196], tmp6964[195], tmp6964[194], tmp6964[193], tmp6964[192], tmp6964[191], tmp6964[190], tmp6964[189], tmp6964[188], tmp6964[187], tmp6964[186], tmp6964[185], tmp6964[184], tmp6964[183], tmp6964[182], tmp6964[181], tmp6964[180], tmp6964[179], tmp6964[178], tmp6964[177], tmp6964[176], tmp6964[175], tmp6964[174], tmp6964[173], tmp6964[172], tmp6964[171], tmp6964[170], tmp6964[169], tmp6964[168], tmp6964[167], tmp6964[166], tmp6964[165], tmp6964[164], tmp6964[163], tmp6964[162], tmp6964[161], tmp6964[160], tmp6964[159], tmp6964[158], tmp6964[157], tmp6964[156], tmp6964[155], tmp6964[154], tmp6964[153], tmp6964[152], tmp6964[151], tmp6964[150], tmp6964[149], tmp6964[148], tmp6964[147], tmp6964[146], tmp6964[145], tmp6964[144], tmp6964[143], tmp6964[142], tmp6964[141], tmp6964[140], tmp6964[139], tmp6964[138], tmp6964[137], tmp6964[136], tmp6964[135], tmp6964[134], tmp6964[133], tmp6964[132], tmp6964[131], tmp6964[130], tmp6964[129], tmp6964[128], tmp6964[127], tmp6964[126], tmp6964[125], tmp6964[124], tmp6964[123], tmp6964[122], tmp6964[121], tmp6964[120], tmp6964[119], tmp6964[118], tmp6964[117], tmp6964[116], tmp6964[115], tmp6964[114], tmp6964[113], tmp6964[112], tmp6964[111], tmp6964[110], tmp6964[109], tmp6964[108], tmp6964[107], tmp6964[106], tmp6964[105], tmp6964[104], tmp6964[103], tmp6964[102], tmp6964[101], tmp6964[100], tmp6964[99], tmp6964[98], tmp6964[97], tmp6964[96], tmp6964[95], tmp6964[94], tmp6964[93], tmp6964[92], tmp6964[91], tmp6964[90], tmp6964[89], tmp6964[88], tmp6964[87], tmp6964[86], tmp6964[85], tmp6964[84], tmp6964[83], tmp6964[82], tmp6964[81], tmp6964[80], tmp6964[79], tmp6964[78], tmp6964[77], tmp6964[76], tmp6964[75], tmp6964[74], tmp6964[73], tmp6964[72], tmp6964[71], tmp6964[70], tmp6964[69], tmp6964[68], tmp6964[67], tmp6964[66], tmp6964[65], tmp6964[64], tmp6964[63], tmp6964[62], tmp6964[61], tmp6964[60], tmp6964[59], tmp6964[58], tmp6964[57], tmp6964[56], tmp6964[55], tmp6964[54], tmp6964[53], tmp6964[52], tmp6964[51], tmp6964[50], tmp6964[49], tmp6964[48], tmp6964[47], tmp6964[46], tmp6964[45], tmp6964[44], tmp6964[43], tmp6964[42], tmp6964[41], tmp6964[40], tmp6964[39], tmp6964[38], tmp6964[37], tmp6964[36], tmp6964[35], tmp6964[34], tmp6964[33], tmp6964[32], tmp6964[31], tmp6964[30], tmp6964[29], tmp6964[28], tmp6964[27], tmp6964[26], tmp6964[25], tmp6964[24], tmp6964[23], tmp6964[22], tmp6964[21], tmp6964[20], tmp6964[19], tmp6964[18], tmp6964[17], tmp6964[16], tmp6964[15], tmp6964[14], tmp6964[13], tmp6964[12], tmp6964[11], tmp6964[10], tmp6964[9], tmp6964[8], tmp6964[7], tmp6964[6], tmp6964[5], tmp6964[4], tmp6964[3], tmp6964[2], tmp6964[1]};
    assign tmp6966 = {tmp6965[255]};
    assign tmp6967 = {tmp6966};
    assign tmp6968 = {tmp6967, tmp6965};
    assign tmp6969 = {tmp18[255]};
    assign tmp6970 = {const_682_0};
    assign tmp6971 = {tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970, tmp6970};
    assign tmp6972 = {tmp6971, const_682_0};
    assign tmp6973 = tmp18 - tmp6972;
    assign tmp6974 = {tmp6973[256]};
    assign tmp6975 = {tmp18[255]};
    assign tmp6976 = ~tmp6975;
    assign tmp6977 = tmp6974 ^ tmp6976;
    assign tmp6978 = {tmp6972[255]};
    assign tmp6979 = ~tmp6978;
    assign tmp6980 = tmp6977 ^ tmp6979;
    assign tmp6981 = tmp18 == _ver_out_tmp_47;
    assign tmp6982 = {const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0, const_685_0};
    assign tmp6983 = {tmp6982, const_684_0};
    assign tmp6984 = tmp6983 - tmp18;
    assign tmp6985 = {const_687_0, const_687_0};
    assign tmp6986 = {tmp6985, const_686_57896044618658097711785492504343953926634992332820282019728792003956564819967};
    assign tmp6987 = tmp6981 ? tmp6986 : tmp6984;
    assign tmp6988 = {const_688_0};
    assign tmp6989 = {tmp6988, tmp18};
    assign tmp6990 = tmp6980 ? tmp6989 : tmp6987;
    assign tmp6991 = {tmp6968[256]};
    assign tmp6992 = {tmp6990[256]};
    assign tmp6993 = tmp6990 - tmp6968;
    assign tmp6994 = {tmp6993[257]};
    assign tmp6995 = {tmp6968[256]};
    assign tmp6996 = ~tmp6995;
    assign tmp6997 = tmp6994 ^ tmp6996;
    assign tmp6998 = {tmp6990[256]};
    assign tmp6999 = ~tmp6998;
    assign tmp7000 = tmp6997 ^ tmp6999;
    assign tmp7001 = tmp6968 == tmp6990;
    assign tmp7002 = tmp7000 | tmp7001;
    assign tmp7003 = tmp6942 & tmp7002;
    assign tmp7004 = ~tmp35;
    assign tmp7005 = ~tmp36;
    assign tmp7006 = tmp7004 & tmp7005;
    assign tmp7007 = ~tmp57;
    assign tmp7008 = tmp7006 & tmp7007;
    assign tmp7009 = ~tmp1034;
    assign tmp7010 = tmp7008 & tmp7009;
    assign tmp7011 = tmp7010 & tmp2071;
    assign tmp7012 = ~tmp2583;
    assign tmp7013 = tmp7011 & tmp7012;
    assign tmp7014 = ~tmp23;
    assign tmp7015 = tmp7013 & tmp7014;
    assign tmp7016 = tmp7015 & cfg_speculative_egest;
    assign tmp7017 = ~tmp6619;
    assign tmp7018 = tmp7016 & tmp7017;
    assign tmp7019 = tmp7018 & tmp7003;
    assign tmp7020 = ~tmp35;
    assign tmp7021 = ~tmp36;
    assign tmp7022 = tmp7020 & tmp7021;
    assign tmp7023 = ~tmp57;
    assign tmp7024 = tmp7022 & tmp7023;
    assign tmp7025 = ~tmp1034;
    assign tmp7026 = tmp7024 & tmp7025;
    assign tmp7027 = tmp7026 & tmp2071;
    assign tmp7028 = ~tmp2583;
    assign tmp7029 = tmp7027 & tmp7028;
    assign tmp7030 = ~tmp23;
    assign tmp7031 = tmp7029 & tmp7030;
    assign tmp7032 = tmp7031 & cfg_speculative_egest;
    assign tmp7033 = ~tmp6619;
    assign tmp7034 = tmp7032 & tmp7033;
    assign tmp7035 = tmp7034 & tmp7003;
    assign tmp7036 = {tmp11[255], tmp11[254], tmp11[253], tmp11[252], tmp11[251], tmp11[250], tmp11[249], tmp11[248], tmp11[247], tmp11[246], tmp11[245], tmp11[244], tmp11[243], tmp11[242], tmp11[241], tmp11[240], tmp11[239], tmp11[238], tmp11[237], tmp11[236], tmp11[235], tmp11[234], tmp11[233], tmp11[232], tmp11[231], tmp11[230], tmp11[229], tmp11[228], tmp11[227], tmp11[226], tmp11[225], tmp11[224], tmp11[223], tmp11[222], tmp11[221], tmp11[220], tmp11[219], tmp11[218], tmp11[217], tmp11[216], tmp11[215], tmp11[214], tmp11[213], tmp11[212], tmp11[211], tmp11[210], tmp11[209], tmp11[208], tmp11[207], tmp11[206], tmp11[205], tmp11[204], tmp11[203], tmp11[202], tmp11[201], tmp11[200], tmp11[199], tmp11[198], tmp11[197], tmp11[196], tmp11[195], tmp11[194], tmp11[193], tmp11[192], tmp11[191], tmp11[190], tmp11[189], tmp11[188], tmp11[187], tmp11[186], tmp11[185], tmp11[184], tmp11[183], tmp11[182], tmp11[181], tmp11[180], tmp11[179], tmp11[178], tmp11[177], tmp11[176], tmp11[175], tmp11[174], tmp11[173], tmp11[172], tmp11[171], tmp11[170], tmp11[169], tmp11[168], tmp11[167], tmp11[166], tmp11[165], tmp11[164], tmp11[163], tmp11[162], tmp11[161], tmp11[160], tmp11[159], tmp11[158], tmp11[157], tmp11[156], tmp11[155], tmp11[154], tmp11[153], tmp11[152], tmp11[151], tmp11[150], tmp11[149], tmp11[148], tmp11[147], tmp11[146], tmp11[145], tmp11[144], tmp11[143], tmp11[142], tmp11[141], tmp11[140], tmp11[139], tmp11[138], tmp11[137], tmp11[136], tmp11[135], tmp11[134], tmp11[133], tmp11[132], tmp11[131], tmp11[130], tmp11[129], tmp11[128], tmp11[127], tmp11[126], tmp11[125], tmp11[124], tmp11[123], tmp11[122], tmp11[121], tmp11[120], tmp11[119], tmp11[118], tmp11[117], tmp11[116], tmp11[115], tmp11[114], tmp11[113], tmp11[112], tmp11[111], tmp11[110], tmp11[109], tmp11[108], tmp11[107], tmp11[106], tmp11[105], tmp11[104], tmp11[103], tmp11[102], tmp11[101], tmp11[100], tmp11[99], tmp11[98], tmp11[97], tmp11[96], tmp11[95], tmp11[94], tmp11[93], tmp11[92], tmp11[91], tmp11[90], tmp11[89], tmp11[88], tmp11[87], tmp11[86], tmp11[85], tmp11[84], tmp11[83], tmp11[82], tmp11[81], tmp11[80], tmp11[79], tmp11[78], tmp11[77], tmp11[76], tmp11[75], tmp11[74], tmp11[73], tmp11[72], tmp11[71], tmp11[70], tmp11[69], tmp11[68], tmp11[67], tmp11[66], tmp11[65], tmp11[64], tmp11[63], tmp11[62], tmp11[61], tmp11[60], tmp11[59], tmp11[58], tmp11[57], tmp11[56], tmp11[55], tmp11[54], tmp11[53], tmp11[52], tmp11[51], tmp11[50], tmp11[49], tmp11[48], tmp11[47], tmp11[46], tmp11[45], tmp11[44], tmp11[43], tmp11[42], tmp11[41], tmp11[40], tmp11[39], tmp11[38], tmp11[37], tmp11[36], tmp11[35], tmp11[34], tmp11[33], tmp11[32], tmp11[31], tmp11[30], tmp11[29], tmp11[28], tmp11[27], tmp11[26], tmp11[25], tmp11[24], tmp11[23], tmp11[22], tmp11[21], tmp11[20], tmp11[19], tmp11[18], tmp11[17], tmp11[16], tmp11[15], tmp11[14], tmp11[13], tmp11[12], tmp11[11], tmp11[10], tmp11[9], tmp11[8], tmp11[7], tmp11[6], tmp11[5], tmp11[4], tmp11[3], tmp11[2], tmp11[1]};
    assign tmp7037 = {tmp7036[254]};
    assign tmp7038 = {tmp7037};
    assign tmp7039 = {tmp7038, tmp7036};
    assign tmp7040 = ~tmp35;
    assign tmp7041 = ~tmp36;
    assign tmp7042 = tmp7040 & tmp7041;
    assign tmp7043 = ~tmp57;
    assign tmp7044 = tmp7042 & tmp7043;
    assign tmp7045 = ~tmp1034;
    assign tmp7046 = tmp7044 & tmp7045;
    assign tmp7047 = tmp7046 & tmp2071;
    assign tmp7048 = ~tmp2583;
    assign tmp7049 = tmp7047 & tmp7048;
    assign tmp7050 = ~tmp23;
    assign tmp7051 = tmp7049 & tmp7050;
    assign tmp7052 = tmp7051 & cfg_speculative_egest;
    assign tmp7053 = ~tmp6619;
    assign tmp7054 = tmp7052 & tmp7053;
    assign tmp7055 = tmp7054 & tmp7003;
    assign tmp7056 = tmp7055 & tmp24;
    assign tmp7057 = {tmp12[255], tmp12[254], tmp12[253], tmp12[252], tmp12[251], tmp12[250], tmp12[249], tmp12[248], tmp12[247], tmp12[246], tmp12[245], tmp12[244], tmp12[243], tmp12[242], tmp12[241], tmp12[240], tmp12[239], tmp12[238], tmp12[237], tmp12[236], tmp12[235], tmp12[234], tmp12[233], tmp12[232], tmp12[231], tmp12[230], tmp12[229], tmp12[228], tmp12[227], tmp12[226], tmp12[225], tmp12[224], tmp12[223], tmp12[222], tmp12[221], tmp12[220], tmp12[219], tmp12[218], tmp12[217], tmp12[216], tmp12[215], tmp12[214], tmp12[213], tmp12[212], tmp12[211], tmp12[210], tmp12[209], tmp12[208], tmp12[207], tmp12[206], tmp12[205], tmp12[204], tmp12[203], tmp12[202], tmp12[201], tmp12[200], tmp12[199], tmp12[198], tmp12[197], tmp12[196], tmp12[195], tmp12[194], tmp12[193], tmp12[192], tmp12[191], tmp12[190], tmp12[189], tmp12[188], tmp12[187], tmp12[186], tmp12[185], tmp12[184], tmp12[183], tmp12[182], tmp12[181], tmp12[180], tmp12[179], tmp12[178], tmp12[177], tmp12[176], tmp12[175], tmp12[174], tmp12[173], tmp12[172], tmp12[171], tmp12[170], tmp12[169], tmp12[168], tmp12[167], tmp12[166], tmp12[165], tmp12[164], tmp12[163], tmp12[162], tmp12[161], tmp12[160], tmp12[159], tmp12[158], tmp12[157], tmp12[156], tmp12[155], tmp12[154], tmp12[153], tmp12[152], tmp12[151], tmp12[150], tmp12[149], tmp12[148], tmp12[147], tmp12[146], tmp12[145], tmp12[144], tmp12[143], tmp12[142], tmp12[141], tmp12[140], tmp12[139], tmp12[138], tmp12[137], tmp12[136], tmp12[135], tmp12[134], tmp12[133], tmp12[132], tmp12[131], tmp12[130], tmp12[129], tmp12[128], tmp12[127], tmp12[126], tmp12[125], tmp12[124], tmp12[123], tmp12[122], tmp12[121], tmp12[120], tmp12[119], tmp12[118], tmp12[117], tmp12[116], tmp12[115], tmp12[114], tmp12[113], tmp12[112], tmp12[111], tmp12[110], tmp12[109], tmp12[108], tmp12[107], tmp12[106], tmp12[105], tmp12[104], tmp12[103], tmp12[102], tmp12[101], tmp12[100], tmp12[99], tmp12[98], tmp12[97], tmp12[96], tmp12[95], tmp12[94], tmp12[93], tmp12[92], tmp12[91], tmp12[90], tmp12[89], tmp12[88], tmp12[87], tmp12[86], tmp12[85], tmp12[84], tmp12[83], tmp12[82], tmp12[81], tmp12[80], tmp12[79], tmp12[78], tmp12[77], tmp12[76], tmp12[75], tmp12[74], tmp12[73], tmp12[72], tmp12[71], tmp12[70], tmp12[69], tmp12[68], tmp12[67], tmp12[66], tmp12[65], tmp12[64], tmp12[63], tmp12[62], tmp12[61], tmp12[60], tmp12[59], tmp12[58], tmp12[57], tmp12[56], tmp12[55], tmp12[54], tmp12[53], tmp12[52], tmp12[51], tmp12[50], tmp12[49], tmp12[48], tmp12[47], tmp12[46], tmp12[45], tmp12[44], tmp12[43], tmp12[42], tmp12[41], tmp12[40], tmp12[39], tmp12[38], tmp12[37], tmp12[36], tmp12[35], tmp12[34], tmp12[33], tmp12[32], tmp12[31], tmp12[30], tmp12[29], tmp12[28], tmp12[27], tmp12[26], tmp12[25], tmp12[24], tmp12[23], tmp12[22], tmp12[21], tmp12[20], tmp12[19], tmp12[18], tmp12[17], tmp12[16], tmp12[15], tmp12[14], tmp12[13], tmp12[12], tmp12[11], tmp12[10], tmp12[9], tmp12[8], tmp12[7], tmp12[6], tmp12[5], tmp12[4], tmp12[3], tmp12[2], tmp12[1]};
    assign tmp7058 = {tmp7057[254]};
    assign tmp7059 = {tmp7058};
    assign tmp7060 = {tmp7059, tmp7057};
    assign tmp7061 = ~tmp35;
    assign tmp7062 = ~tmp36;
    assign tmp7063 = tmp7061 & tmp7062;
    assign tmp7064 = ~tmp57;
    assign tmp7065 = tmp7063 & tmp7064;
    assign tmp7066 = ~tmp1034;
    assign tmp7067 = tmp7065 & tmp7066;
    assign tmp7068 = tmp7067 & tmp2071;
    assign tmp7069 = ~tmp2583;
    assign tmp7070 = tmp7068 & tmp7069;
    assign tmp7071 = ~tmp23;
    assign tmp7072 = tmp7070 & tmp7071;
    assign tmp7073 = tmp7072 & cfg_speculative_egest;
    assign tmp7074 = ~tmp6619;
    assign tmp7075 = tmp7073 & tmp7074;
    assign tmp7076 = tmp7075 & tmp7003;
    assign tmp7077 = tmp7076 & tmp24;
    assign tmp7078 = {tmp13[255], tmp13[254], tmp13[253], tmp13[252], tmp13[251], tmp13[250], tmp13[249], tmp13[248], tmp13[247], tmp13[246], tmp13[245], tmp13[244], tmp13[243], tmp13[242], tmp13[241], tmp13[240], tmp13[239], tmp13[238], tmp13[237], tmp13[236], tmp13[235], tmp13[234], tmp13[233], tmp13[232], tmp13[231], tmp13[230], tmp13[229], tmp13[228], tmp13[227], tmp13[226], tmp13[225], tmp13[224], tmp13[223], tmp13[222], tmp13[221], tmp13[220], tmp13[219], tmp13[218], tmp13[217], tmp13[216], tmp13[215], tmp13[214], tmp13[213], tmp13[212], tmp13[211], tmp13[210], tmp13[209], tmp13[208], tmp13[207], tmp13[206], tmp13[205], tmp13[204], tmp13[203], tmp13[202], tmp13[201], tmp13[200], tmp13[199], tmp13[198], tmp13[197], tmp13[196], tmp13[195], tmp13[194], tmp13[193], tmp13[192], tmp13[191], tmp13[190], tmp13[189], tmp13[188], tmp13[187], tmp13[186], tmp13[185], tmp13[184], tmp13[183], tmp13[182], tmp13[181], tmp13[180], tmp13[179], tmp13[178], tmp13[177], tmp13[176], tmp13[175], tmp13[174], tmp13[173], tmp13[172], tmp13[171], tmp13[170], tmp13[169], tmp13[168], tmp13[167], tmp13[166], tmp13[165], tmp13[164], tmp13[163], tmp13[162], tmp13[161], tmp13[160], tmp13[159], tmp13[158], tmp13[157], tmp13[156], tmp13[155], tmp13[154], tmp13[153], tmp13[152], tmp13[151], tmp13[150], tmp13[149], tmp13[148], tmp13[147], tmp13[146], tmp13[145], tmp13[144], tmp13[143], tmp13[142], tmp13[141], tmp13[140], tmp13[139], tmp13[138], tmp13[137], tmp13[136], tmp13[135], tmp13[134], tmp13[133], tmp13[132], tmp13[131], tmp13[130], tmp13[129], tmp13[128], tmp13[127], tmp13[126], tmp13[125], tmp13[124], tmp13[123], tmp13[122], tmp13[121], tmp13[120], tmp13[119], tmp13[118], tmp13[117], tmp13[116], tmp13[115], tmp13[114], tmp13[113], tmp13[112], tmp13[111], tmp13[110], tmp13[109], tmp13[108], tmp13[107], tmp13[106], tmp13[105], tmp13[104], tmp13[103], tmp13[102], tmp13[101], tmp13[100], tmp13[99], tmp13[98], tmp13[97], tmp13[96], tmp13[95], tmp13[94], tmp13[93], tmp13[92], tmp13[91], tmp13[90], tmp13[89], tmp13[88], tmp13[87], tmp13[86], tmp13[85], tmp13[84], tmp13[83], tmp13[82], tmp13[81], tmp13[80], tmp13[79], tmp13[78], tmp13[77], tmp13[76], tmp13[75], tmp13[74], tmp13[73], tmp13[72], tmp13[71], tmp13[70], tmp13[69], tmp13[68], tmp13[67], tmp13[66], tmp13[65], tmp13[64], tmp13[63], tmp13[62], tmp13[61], tmp13[60], tmp13[59], tmp13[58], tmp13[57], tmp13[56], tmp13[55], tmp13[54], tmp13[53], tmp13[52], tmp13[51], tmp13[50], tmp13[49], tmp13[48], tmp13[47], tmp13[46], tmp13[45], tmp13[44], tmp13[43], tmp13[42], tmp13[41], tmp13[40], tmp13[39], tmp13[38], tmp13[37], tmp13[36], tmp13[35], tmp13[34], tmp13[33], tmp13[32], tmp13[31], tmp13[30], tmp13[29], tmp13[28], tmp13[27], tmp13[26], tmp13[25], tmp13[24], tmp13[23], tmp13[22], tmp13[21], tmp13[20], tmp13[19], tmp13[18], tmp13[17], tmp13[16], tmp13[15], tmp13[14], tmp13[13], tmp13[12], tmp13[11], tmp13[10], tmp13[9], tmp13[8], tmp13[7], tmp13[6], tmp13[5], tmp13[4], tmp13[3], tmp13[2], tmp13[1]};
    assign tmp7079 = {tmp7078[254]};
    assign tmp7080 = {tmp7079};
    assign tmp7081 = {tmp7080, tmp7078};
    assign tmp7082 = ~tmp35;
    assign tmp7083 = ~tmp36;
    assign tmp7084 = tmp7082 & tmp7083;
    assign tmp7085 = ~tmp57;
    assign tmp7086 = tmp7084 & tmp7085;
    assign tmp7087 = ~tmp1034;
    assign tmp7088 = tmp7086 & tmp7087;
    assign tmp7089 = tmp7088 & tmp2071;
    assign tmp7090 = ~tmp2583;
    assign tmp7091 = tmp7089 & tmp7090;
    assign tmp7092 = ~tmp23;
    assign tmp7093 = tmp7091 & tmp7092;
    assign tmp7094 = tmp7093 & cfg_speculative_egest;
    assign tmp7095 = ~tmp6619;
    assign tmp7096 = tmp7094 & tmp7095;
    assign tmp7097 = tmp7096 & tmp7003;
    assign tmp7098 = tmp7097 & tmp24;
    assign tmp7099 = {tmp14[255], tmp14[254], tmp14[253], tmp14[252], tmp14[251], tmp14[250], tmp14[249], tmp14[248], tmp14[247], tmp14[246], tmp14[245], tmp14[244], tmp14[243], tmp14[242], tmp14[241], tmp14[240], tmp14[239], tmp14[238], tmp14[237], tmp14[236], tmp14[235], tmp14[234], tmp14[233], tmp14[232], tmp14[231], tmp14[230], tmp14[229], tmp14[228], tmp14[227], tmp14[226], tmp14[225], tmp14[224], tmp14[223], tmp14[222], tmp14[221], tmp14[220], tmp14[219], tmp14[218], tmp14[217], tmp14[216], tmp14[215], tmp14[214], tmp14[213], tmp14[212], tmp14[211], tmp14[210], tmp14[209], tmp14[208], tmp14[207], tmp14[206], tmp14[205], tmp14[204], tmp14[203], tmp14[202], tmp14[201], tmp14[200], tmp14[199], tmp14[198], tmp14[197], tmp14[196], tmp14[195], tmp14[194], tmp14[193], tmp14[192], tmp14[191], tmp14[190], tmp14[189], tmp14[188], tmp14[187], tmp14[186], tmp14[185], tmp14[184], tmp14[183], tmp14[182], tmp14[181], tmp14[180], tmp14[179], tmp14[178], tmp14[177], tmp14[176], tmp14[175], tmp14[174], tmp14[173], tmp14[172], tmp14[171], tmp14[170], tmp14[169], tmp14[168], tmp14[167], tmp14[166], tmp14[165], tmp14[164], tmp14[163], tmp14[162], tmp14[161], tmp14[160], tmp14[159], tmp14[158], tmp14[157], tmp14[156], tmp14[155], tmp14[154], tmp14[153], tmp14[152], tmp14[151], tmp14[150], tmp14[149], tmp14[148], tmp14[147], tmp14[146], tmp14[145], tmp14[144], tmp14[143], tmp14[142], tmp14[141], tmp14[140], tmp14[139], tmp14[138], tmp14[137], tmp14[136], tmp14[135], tmp14[134], tmp14[133], tmp14[132], tmp14[131], tmp14[130], tmp14[129], tmp14[128], tmp14[127], tmp14[126], tmp14[125], tmp14[124], tmp14[123], tmp14[122], tmp14[121], tmp14[120], tmp14[119], tmp14[118], tmp14[117], tmp14[116], tmp14[115], tmp14[114], tmp14[113], tmp14[112], tmp14[111], tmp14[110], tmp14[109], tmp14[108], tmp14[107], tmp14[106], tmp14[105], tmp14[104], tmp14[103], tmp14[102], tmp14[101], tmp14[100], tmp14[99], tmp14[98], tmp14[97], tmp14[96], tmp14[95], tmp14[94], tmp14[93], tmp14[92], tmp14[91], tmp14[90], tmp14[89], tmp14[88], tmp14[87], tmp14[86], tmp14[85], tmp14[84], tmp14[83], tmp14[82], tmp14[81], tmp14[80], tmp14[79], tmp14[78], tmp14[77], tmp14[76], tmp14[75], tmp14[74], tmp14[73], tmp14[72], tmp14[71], tmp14[70], tmp14[69], tmp14[68], tmp14[67], tmp14[66], tmp14[65], tmp14[64], tmp14[63], tmp14[62], tmp14[61], tmp14[60], tmp14[59], tmp14[58], tmp14[57], tmp14[56], tmp14[55], tmp14[54], tmp14[53], tmp14[52], tmp14[51], tmp14[50], tmp14[49], tmp14[48], tmp14[47], tmp14[46], tmp14[45], tmp14[44], tmp14[43], tmp14[42], tmp14[41], tmp14[40], tmp14[39], tmp14[38], tmp14[37], tmp14[36], tmp14[35], tmp14[34], tmp14[33], tmp14[32], tmp14[31], tmp14[30], tmp14[29], tmp14[28], tmp14[27], tmp14[26], tmp14[25], tmp14[24], tmp14[23], tmp14[22], tmp14[21], tmp14[20], tmp14[19], tmp14[18], tmp14[17], tmp14[16], tmp14[15], tmp14[14], tmp14[13], tmp14[12], tmp14[11], tmp14[10], tmp14[9], tmp14[8], tmp14[7], tmp14[6], tmp14[5], tmp14[4], tmp14[3], tmp14[2], tmp14[1]};
    assign tmp7100 = {tmp7099[254]};
    assign tmp7101 = {tmp7100};
    assign tmp7102 = {tmp7101, tmp7099};
    assign tmp7103 = ~tmp35;
    assign tmp7104 = ~tmp36;
    assign tmp7105 = tmp7103 & tmp7104;
    assign tmp7106 = ~tmp57;
    assign tmp7107 = tmp7105 & tmp7106;
    assign tmp7108 = ~tmp1034;
    assign tmp7109 = tmp7107 & tmp7108;
    assign tmp7110 = tmp7109 & tmp2071;
    assign tmp7111 = ~tmp2583;
    assign tmp7112 = tmp7110 & tmp7111;
    assign tmp7113 = ~tmp23;
    assign tmp7114 = tmp7112 & tmp7113;
    assign tmp7115 = tmp7114 & cfg_speculative_egest;
    assign tmp7116 = ~tmp6619;
    assign tmp7117 = tmp7115 & tmp7116;
    assign tmp7118 = tmp7117 & tmp7003;
    assign tmp7119 = tmp7118 & tmp24;
    assign tmp7120 = {tmp15[254], tmp15[253], tmp15[252], tmp15[251], tmp15[250], tmp15[249], tmp15[248], tmp15[247], tmp15[246], tmp15[245], tmp15[244], tmp15[243], tmp15[242], tmp15[241], tmp15[240], tmp15[239], tmp15[238], tmp15[237], tmp15[236], tmp15[235], tmp15[234], tmp15[233], tmp15[232], tmp15[231], tmp15[230], tmp15[229], tmp15[228], tmp15[227], tmp15[226], tmp15[225], tmp15[224], tmp15[223], tmp15[222], tmp15[221], tmp15[220], tmp15[219], tmp15[218], tmp15[217], tmp15[216], tmp15[215], tmp15[214], tmp15[213], tmp15[212], tmp15[211], tmp15[210], tmp15[209], tmp15[208], tmp15[207], tmp15[206], tmp15[205], tmp15[204], tmp15[203], tmp15[202], tmp15[201], tmp15[200], tmp15[199], tmp15[198], tmp15[197], tmp15[196], tmp15[195], tmp15[194], tmp15[193], tmp15[192], tmp15[191], tmp15[190], tmp15[189], tmp15[188], tmp15[187], tmp15[186], tmp15[185], tmp15[184], tmp15[183], tmp15[182], tmp15[181], tmp15[180], tmp15[179], tmp15[178], tmp15[177], tmp15[176], tmp15[175], tmp15[174], tmp15[173], tmp15[172], tmp15[171], tmp15[170], tmp15[169], tmp15[168], tmp15[167], tmp15[166], tmp15[165], tmp15[164], tmp15[163], tmp15[162], tmp15[161], tmp15[160], tmp15[159], tmp15[158], tmp15[157], tmp15[156], tmp15[155], tmp15[154], tmp15[153], tmp15[152], tmp15[151], tmp15[150], tmp15[149], tmp15[148], tmp15[147], tmp15[146], tmp15[145], tmp15[144], tmp15[143], tmp15[142], tmp15[141], tmp15[140], tmp15[139], tmp15[138], tmp15[137], tmp15[136], tmp15[135], tmp15[134], tmp15[133], tmp15[132], tmp15[131], tmp15[130], tmp15[129], tmp15[128], tmp15[127], tmp15[126], tmp15[125], tmp15[124], tmp15[123], tmp15[122], tmp15[121], tmp15[120], tmp15[119], tmp15[118], tmp15[117], tmp15[116], tmp15[115], tmp15[114], tmp15[113], tmp15[112], tmp15[111], tmp15[110], tmp15[109], tmp15[108], tmp15[107], tmp15[106], tmp15[105], tmp15[104], tmp15[103], tmp15[102], tmp15[101], tmp15[100], tmp15[99], tmp15[98], tmp15[97], tmp15[96], tmp15[95], tmp15[94], tmp15[93], tmp15[92], tmp15[91], tmp15[90], tmp15[89], tmp15[88], tmp15[87], tmp15[86], tmp15[85], tmp15[84], tmp15[83], tmp15[82], tmp15[81], tmp15[80], tmp15[79], tmp15[78], tmp15[77], tmp15[76], tmp15[75], tmp15[74], tmp15[73], tmp15[72], tmp15[71], tmp15[70], tmp15[69], tmp15[68], tmp15[67], tmp15[66], tmp15[65], tmp15[64], tmp15[63], tmp15[62], tmp15[61], tmp15[60], tmp15[59], tmp15[58], tmp15[57], tmp15[56], tmp15[55], tmp15[54], tmp15[53], tmp15[52], tmp15[51], tmp15[50], tmp15[49], tmp15[48], tmp15[47], tmp15[46], tmp15[45], tmp15[44], tmp15[43], tmp15[42], tmp15[41], tmp15[40], tmp15[39], tmp15[38], tmp15[37], tmp15[36], tmp15[35], tmp15[34], tmp15[33], tmp15[32], tmp15[31], tmp15[30], tmp15[29], tmp15[28], tmp15[27], tmp15[26], tmp15[25], tmp15[24], tmp15[23], tmp15[22], tmp15[21], tmp15[20], tmp15[19], tmp15[18], tmp15[17], tmp15[16], tmp15[15], tmp15[14], tmp15[13], tmp15[12], tmp15[11], tmp15[10], tmp15[9], tmp15[8], tmp15[7], tmp15[6], tmp15[5], tmp15[4], tmp15[3], tmp15[2], tmp15[1], tmp15[0]};
    assign tmp7121 = {tmp7120, const_691_0};
    assign tmp7122 = {const_692_0};
    assign tmp7123 = {tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122, tmp7122};
    assign tmp7124 = {tmp7123, const_692_0};
    assign tmp7125 = {tmp15[255]};
    assign tmp7126 = tmp7124 - tmp15;
    assign tmp7127 = {tmp7126[256]};
    assign tmp7128 = {tmp7124[255]};
    assign tmp7129 = ~tmp7128;
    assign tmp7130 = tmp7127 ^ tmp7129;
    assign tmp7131 = {tmp15[255]};
    assign tmp7132 = ~tmp7131;
    assign tmp7133 = tmp7130 ^ tmp7132;
    assign tmp7134 = {tmp7121[255]};
    assign tmp7135 = {const_693_0};
    assign tmp7136 = {tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135, tmp7135};
    assign tmp7137 = {tmp7136, const_693_0};
    assign tmp7138 = tmp7121 - tmp7137;
    assign tmp7139 = {tmp7138[256]};
    assign tmp7140 = {tmp7121[255]};
    assign tmp7141 = ~tmp7140;
    assign tmp7142 = tmp7139 ^ tmp7141;
    assign tmp7143 = {tmp7137[255]};
    assign tmp7144 = ~tmp7143;
    assign tmp7145 = tmp7142 ^ tmp7144;
    assign tmp7146 = tmp7133 & tmp7145;
    assign tmp7147 = {tmp15[255]};
    assign tmp7148 = {const_694_0};
    assign tmp7149 = {tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148, tmp7148};
    assign tmp7150 = {tmp7149, const_694_0};
    assign tmp7151 = tmp15 - tmp7150;
    assign tmp7152 = {tmp7151[256]};
    assign tmp7153 = {tmp15[255]};
    assign tmp7154 = ~tmp7153;
    assign tmp7155 = tmp7152 ^ tmp7154;
    assign tmp7156 = {tmp7150[255]};
    assign tmp7157 = ~tmp7156;
    assign tmp7158 = tmp7155 ^ tmp7157;
    assign tmp7159 = {const_695_0};
    assign tmp7160 = {tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159, tmp7159};
    assign tmp7161 = {tmp7160, const_695_0};
    assign tmp7162 = {tmp7121[255]};
    assign tmp7163 = tmp7161 - tmp7121;
    assign tmp7164 = {tmp7163[256]};
    assign tmp7165 = {tmp7161[255]};
    assign tmp7166 = ~tmp7165;
    assign tmp7167 = tmp7164 ^ tmp7166;
    assign tmp7168 = {tmp7121[255]};
    assign tmp7169 = ~tmp7168;
    assign tmp7170 = tmp7167 ^ tmp7169;
    assign tmp7171 = tmp7161 == tmp7121;
    assign tmp7172 = tmp7170 | tmp7171;
    assign tmp7173 = tmp7158 & tmp7172;
    assign tmp7174 = tmp7146 ? const_696_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp7121;
    assign tmp7175 = tmp7173 ? _ver_out_tmp_54 : tmp7174;
    assign tmp7176 = ~tmp35;
    assign tmp7177 = ~tmp36;
    assign tmp7178 = tmp7176 & tmp7177;
    assign tmp7179 = ~tmp57;
    assign tmp7180 = tmp7178 & tmp7179;
    assign tmp7181 = ~tmp1034;
    assign tmp7182 = tmp7180 & tmp7181;
    assign tmp7183 = tmp7182 & tmp2071;
    assign tmp7184 = ~tmp2583;
    assign tmp7185 = tmp7183 & tmp7184;
    assign tmp7186 = ~tmp23;
    assign tmp7187 = tmp7185 & tmp7186;
    assign tmp7188 = tmp7187 & cfg_speculative_egest;
    assign tmp7189 = ~tmp6619;
    assign tmp7190 = tmp7188 & tmp7189;
    assign tmp7191 = tmp7190 & tmp7003;
    assign tmp7192 = ~tmp24;
    assign tmp7193 = tmp7191 & tmp7192;
    assign tmp7194 = {tmp16[254], tmp16[253], tmp16[252], tmp16[251], tmp16[250], tmp16[249], tmp16[248], tmp16[247], tmp16[246], tmp16[245], tmp16[244], tmp16[243], tmp16[242], tmp16[241], tmp16[240], tmp16[239], tmp16[238], tmp16[237], tmp16[236], tmp16[235], tmp16[234], tmp16[233], tmp16[232], tmp16[231], tmp16[230], tmp16[229], tmp16[228], tmp16[227], tmp16[226], tmp16[225], tmp16[224], tmp16[223], tmp16[222], tmp16[221], tmp16[220], tmp16[219], tmp16[218], tmp16[217], tmp16[216], tmp16[215], tmp16[214], tmp16[213], tmp16[212], tmp16[211], tmp16[210], tmp16[209], tmp16[208], tmp16[207], tmp16[206], tmp16[205], tmp16[204], tmp16[203], tmp16[202], tmp16[201], tmp16[200], tmp16[199], tmp16[198], tmp16[197], tmp16[196], tmp16[195], tmp16[194], tmp16[193], tmp16[192], tmp16[191], tmp16[190], tmp16[189], tmp16[188], tmp16[187], tmp16[186], tmp16[185], tmp16[184], tmp16[183], tmp16[182], tmp16[181], tmp16[180], tmp16[179], tmp16[178], tmp16[177], tmp16[176], tmp16[175], tmp16[174], tmp16[173], tmp16[172], tmp16[171], tmp16[170], tmp16[169], tmp16[168], tmp16[167], tmp16[166], tmp16[165], tmp16[164], tmp16[163], tmp16[162], tmp16[161], tmp16[160], tmp16[159], tmp16[158], tmp16[157], tmp16[156], tmp16[155], tmp16[154], tmp16[153], tmp16[152], tmp16[151], tmp16[150], tmp16[149], tmp16[148], tmp16[147], tmp16[146], tmp16[145], tmp16[144], tmp16[143], tmp16[142], tmp16[141], tmp16[140], tmp16[139], tmp16[138], tmp16[137], tmp16[136], tmp16[135], tmp16[134], tmp16[133], tmp16[132], tmp16[131], tmp16[130], tmp16[129], tmp16[128], tmp16[127], tmp16[126], tmp16[125], tmp16[124], tmp16[123], tmp16[122], tmp16[121], tmp16[120], tmp16[119], tmp16[118], tmp16[117], tmp16[116], tmp16[115], tmp16[114], tmp16[113], tmp16[112], tmp16[111], tmp16[110], tmp16[109], tmp16[108], tmp16[107], tmp16[106], tmp16[105], tmp16[104], tmp16[103], tmp16[102], tmp16[101], tmp16[100], tmp16[99], tmp16[98], tmp16[97], tmp16[96], tmp16[95], tmp16[94], tmp16[93], tmp16[92], tmp16[91], tmp16[90], tmp16[89], tmp16[88], tmp16[87], tmp16[86], tmp16[85], tmp16[84], tmp16[83], tmp16[82], tmp16[81], tmp16[80], tmp16[79], tmp16[78], tmp16[77], tmp16[76], tmp16[75], tmp16[74], tmp16[73], tmp16[72], tmp16[71], tmp16[70], tmp16[69], tmp16[68], tmp16[67], tmp16[66], tmp16[65], tmp16[64], tmp16[63], tmp16[62], tmp16[61], tmp16[60], tmp16[59], tmp16[58], tmp16[57], tmp16[56], tmp16[55], tmp16[54], tmp16[53], tmp16[52], tmp16[51], tmp16[50], tmp16[49], tmp16[48], tmp16[47], tmp16[46], tmp16[45], tmp16[44], tmp16[43], tmp16[42], tmp16[41], tmp16[40], tmp16[39], tmp16[38], tmp16[37], tmp16[36], tmp16[35], tmp16[34], tmp16[33], tmp16[32], tmp16[31], tmp16[30], tmp16[29], tmp16[28], tmp16[27], tmp16[26], tmp16[25], tmp16[24], tmp16[23], tmp16[22], tmp16[21], tmp16[20], tmp16[19], tmp16[18], tmp16[17], tmp16[16], tmp16[15], tmp16[14], tmp16[13], tmp16[12], tmp16[11], tmp16[10], tmp16[9], tmp16[8], tmp16[7], tmp16[6], tmp16[5], tmp16[4], tmp16[3], tmp16[2], tmp16[1], tmp16[0]};
    assign tmp7195 = {tmp7194, const_698_0};
    assign tmp7196 = {const_699_0};
    assign tmp7197 = {tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196, tmp7196};
    assign tmp7198 = {tmp7197, const_699_0};
    assign tmp7199 = {tmp16[255]};
    assign tmp7200 = tmp7198 - tmp16;
    assign tmp7201 = {tmp7200[256]};
    assign tmp7202 = {tmp7198[255]};
    assign tmp7203 = ~tmp7202;
    assign tmp7204 = tmp7201 ^ tmp7203;
    assign tmp7205 = {tmp16[255]};
    assign tmp7206 = ~tmp7205;
    assign tmp7207 = tmp7204 ^ tmp7206;
    assign tmp7208 = {tmp7195[255]};
    assign tmp7209 = {const_700_0};
    assign tmp7210 = {tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209, tmp7209};
    assign tmp7211 = {tmp7210, const_700_0};
    assign tmp7212 = tmp7195 - tmp7211;
    assign tmp7213 = {tmp7212[256]};
    assign tmp7214 = {tmp7195[255]};
    assign tmp7215 = ~tmp7214;
    assign tmp7216 = tmp7213 ^ tmp7215;
    assign tmp7217 = {tmp7211[255]};
    assign tmp7218 = ~tmp7217;
    assign tmp7219 = tmp7216 ^ tmp7218;
    assign tmp7220 = tmp7207 & tmp7219;
    assign tmp7221 = {tmp16[255]};
    assign tmp7222 = {const_701_0};
    assign tmp7223 = {tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222, tmp7222};
    assign tmp7224 = {tmp7223, const_701_0};
    assign tmp7225 = tmp16 - tmp7224;
    assign tmp7226 = {tmp7225[256]};
    assign tmp7227 = {tmp16[255]};
    assign tmp7228 = ~tmp7227;
    assign tmp7229 = tmp7226 ^ tmp7228;
    assign tmp7230 = {tmp7224[255]};
    assign tmp7231 = ~tmp7230;
    assign tmp7232 = tmp7229 ^ tmp7231;
    assign tmp7233 = {const_702_0};
    assign tmp7234 = {tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233, tmp7233};
    assign tmp7235 = {tmp7234, const_702_0};
    assign tmp7236 = {tmp7195[255]};
    assign tmp7237 = tmp7235 - tmp7195;
    assign tmp7238 = {tmp7237[256]};
    assign tmp7239 = {tmp7235[255]};
    assign tmp7240 = ~tmp7239;
    assign tmp7241 = tmp7238 ^ tmp7240;
    assign tmp7242 = {tmp7195[255]};
    assign tmp7243 = ~tmp7242;
    assign tmp7244 = tmp7241 ^ tmp7243;
    assign tmp7245 = tmp7235 == tmp7195;
    assign tmp7246 = tmp7244 | tmp7245;
    assign tmp7247 = tmp7232 & tmp7246;
    assign tmp7248 = tmp7220 ? const_703_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp7195;
    assign tmp7249 = tmp7247 ? _ver_out_tmp_58 : tmp7248;
    assign tmp7250 = ~tmp35;
    assign tmp7251 = ~tmp36;
    assign tmp7252 = tmp7250 & tmp7251;
    assign tmp7253 = ~tmp57;
    assign tmp7254 = tmp7252 & tmp7253;
    assign tmp7255 = ~tmp1034;
    assign tmp7256 = tmp7254 & tmp7255;
    assign tmp7257 = tmp7256 & tmp2071;
    assign tmp7258 = ~tmp2583;
    assign tmp7259 = tmp7257 & tmp7258;
    assign tmp7260 = ~tmp23;
    assign tmp7261 = tmp7259 & tmp7260;
    assign tmp7262 = tmp7261 & cfg_speculative_egest;
    assign tmp7263 = ~tmp6619;
    assign tmp7264 = tmp7262 & tmp7263;
    assign tmp7265 = tmp7264 & tmp7003;
    assign tmp7266 = ~tmp24;
    assign tmp7267 = tmp7265 & tmp7266;
    assign tmp7268 = {tmp17[254], tmp17[253], tmp17[252], tmp17[251], tmp17[250], tmp17[249], tmp17[248], tmp17[247], tmp17[246], tmp17[245], tmp17[244], tmp17[243], tmp17[242], tmp17[241], tmp17[240], tmp17[239], tmp17[238], tmp17[237], tmp17[236], tmp17[235], tmp17[234], tmp17[233], tmp17[232], tmp17[231], tmp17[230], tmp17[229], tmp17[228], tmp17[227], tmp17[226], tmp17[225], tmp17[224], tmp17[223], tmp17[222], tmp17[221], tmp17[220], tmp17[219], tmp17[218], tmp17[217], tmp17[216], tmp17[215], tmp17[214], tmp17[213], tmp17[212], tmp17[211], tmp17[210], tmp17[209], tmp17[208], tmp17[207], tmp17[206], tmp17[205], tmp17[204], tmp17[203], tmp17[202], tmp17[201], tmp17[200], tmp17[199], tmp17[198], tmp17[197], tmp17[196], tmp17[195], tmp17[194], tmp17[193], tmp17[192], tmp17[191], tmp17[190], tmp17[189], tmp17[188], tmp17[187], tmp17[186], tmp17[185], tmp17[184], tmp17[183], tmp17[182], tmp17[181], tmp17[180], tmp17[179], tmp17[178], tmp17[177], tmp17[176], tmp17[175], tmp17[174], tmp17[173], tmp17[172], tmp17[171], tmp17[170], tmp17[169], tmp17[168], tmp17[167], tmp17[166], tmp17[165], tmp17[164], tmp17[163], tmp17[162], tmp17[161], tmp17[160], tmp17[159], tmp17[158], tmp17[157], tmp17[156], tmp17[155], tmp17[154], tmp17[153], tmp17[152], tmp17[151], tmp17[150], tmp17[149], tmp17[148], tmp17[147], tmp17[146], tmp17[145], tmp17[144], tmp17[143], tmp17[142], tmp17[141], tmp17[140], tmp17[139], tmp17[138], tmp17[137], tmp17[136], tmp17[135], tmp17[134], tmp17[133], tmp17[132], tmp17[131], tmp17[130], tmp17[129], tmp17[128], tmp17[127], tmp17[126], tmp17[125], tmp17[124], tmp17[123], tmp17[122], tmp17[121], tmp17[120], tmp17[119], tmp17[118], tmp17[117], tmp17[116], tmp17[115], tmp17[114], tmp17[113], tmp17[112], tmp17[111], tmp17[110], tmp17[109], tmp17[108], tmp17[107], tmp17[106], tmp17[105], tmp17[104], tmp17[103], tmp17[102], tmp17[101], tmp17[100], tmp17[99], tmp17[98], tmp17[97], tmp17[96], tmp17[95], tmp17[94], tmp17[93], tmp17[92], tmp17[91], tmp17[90], tmp17[89], tmp17[88], tmp17[87], tmp17[86], tmp17[85], tmp17[84], tmp17[83], tmp17[82], tmp17[81], tmp17[80], tmp17[79], tmp17[78], tmp17[77], tmp17[76], tmp17[75], tmp17[74], tmp17[73], tmp17[72], tmp17[71], tmp17[70], tmp17[69], tmp17[68], tmp17[67], tmp17[66], tmp17[65], tmp17[64], tmp17[63], tmp17[62], tmp17[61], tmp17[60], tmp17[59], tmp17[58], tmp17[57], tmp17[56], tmp17[55], tmp17[54], tmp17[53], tmp17[52], tmp17[51], tmp17[50], tmp17[49], tmp17[48], tmp17[47], tmp17[46], tmp17[45], tmp17[44], tmp17[43], tmp17[42], tmp17[41], tmp17[40], tmp17[39], tmp17[38], tmp17[37], tmp17[36], tmp17[35], tmp17[34], tmp17[33], tmp17[32], tmp17[31], tmp17[30], tmp17[29], tmp17[28], tmp17[27], tmp17[26], tmp17[25], tmp17[24], tmp17[23], tmp17[22], tmp17[21], tmp17[20], tmp17[19], tmp17[18], tmp17[17], tmp17[16], tmp17[15], tmp17[14], tmp17[13], tmp17[12], tmp17[11], tmp17[10], tmp17[9], tmp17[8], tmp17[7], tmp17[6], tmp17[5], tmp17[4], tmp17[3], tmp17[2], tmp17[1], tmp17[0]};
    assign tmp7269 = {tmp7268, const_705_0};
    assign tmp7270 = {const_706_0};
    assign tmp7271 = {tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270, tmp7270};
    assign tmp7272 = {tmp7271, const_706_0};
    assign tmp7273 = {tmp17[255]};
    assign tmp7274 = tmp7272 - tmp17;
    assign tmp7275 = {tmp7274[256]};
    assign tmp7276 = {tmp7272[255]};
    assign tmp7277 = ~tmp7276;
    assign tmp7278 = tmp7275 ^ tmp7277;
    assign tmp7279 = {tmp17[255]};
    assign tmp7280 = ~tmp7279;
    assign tmp7281 = tmp7278 ^ tmp7280;
    assign tmp7282 = {tmp7269[255]};
    assign tmp7283 = {const_707_0};
    assign tmp7284 = {tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283, tmp7283};
    assign tmp7285 = {tmp7284, const_707_0};
    assign tmp7286 = tmp7269 - tmp7285;
    assign tmp7287 = {tmp7286[256]};
    assign tmp7288 = {tmp7269[255]};
    assign tmp7289 = ~tmp7288;
    assign tmp7290 = tmp7287 ^ tmp7289;
    assign tmp7291 = {tmp7285[255]};
    assign tmp7292 = ~tmp7291;
    assign tmp7293 = tmp7290 ^ tmp7292;
    assign tmp7294 = tmp7281 & tmp7293;
    assign tmp7295 = {tmp17[255]};
    assign tmp7296 = {const_708_0};
    assign tmp7297 = {tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296, tmp7296};
    assign tmp7298 = {tmp7297, const_708_0};
    assign tmp7299 = tmp17 - tmp7298;
    assign tmp7300 = {tmp7299[256]};
    assign tmp7301 = {tmp17[255]};
    assign tmp7302 = ~tmp7301;
    assign tmp7303 = tmp7300 ^ tmp7302;
    assign tmp7304 = {tmp7298[255]};
    assign tmp7305 = ~tmp7304;
    assign tmp7306 = tmp7303 ^ tmp7305;
    assign tmp7307 = {const_709_0};
    assign tmp7308 = {tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307, tmp7307};
    assign tmp7309 = {tmp7308, const_709_0};
    assign tmp7310 = {tmp7269[255]};
    assign tmp7311 = tmp7309 - tmp7269;
    assign tmp7312 = {tmp7311[256]};
    assign tmp7313 = {tmp7309[255]};
    assign tmp7314 = ~tmp7313;
    assign tmp7315 = tmp7312 ^ tmp7314;
    assign tmp7316 = {tmp7269[255]};
    assign tmp7317 = ~tmp7316;
    assign tmp7318 = tmp7315 ^ tmp7317;
    assign tmp7319 = tmp7309 == tmp7269;
    assign tmp7320 = tmp7318 | tmp7319;
    assign tmp7321 = tmp7306 & tmp7320;
    assign tmp7322 = tmp7294 ? const_710_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp7269;
    assign tmp7323 = tmp7321 ? _ver_out_tmp_1 : tmp7322;
    assign tmp7324 = ~tmp35;
    assign tmp7325 = ~tmp36;
    assign tmp7326 = tmp7324 & tmp7325;
    assign tmp7327 = ~tmp57;
    assign tmp7328 = tmp7326 & tmp7327;
    assign tmp7329 = ~tmp1034;
    assign tmp7330 = tmp7328 & tmp7329;
    assign tmp7331 = tmp7330 & tmp2071;
    assign tmp7332 = ~tmp2583;
    assign tmp7333 = tmp7331 & tmp7332;
    assign tmp7334 = ~tmp23;
    assign tmp7335 = tmp7333 & tmp7334;
    assign tmp7336 = tmp7335 & cfg_speculative_egest;
    assign tmp7337 = ~tmp6619;
    assign tmp7338 = tmp7336 & tmp7337;
    assign tmp7339 = tmp7338 & tmp7003;
    assign tmp7340 = ~tmp24;
    assign tmp7341 = tmp7339 & tmp7340;
    assign tmp7342 = {tmp18[254], tmp18[253], tmp18[252], tmp18[251], tmp18[250], tmp18[249], tmp18[248], tmp18[247], tmp18[246], tmp18[245], tmp18[244], tmp18[243], tmp18[242], tmp18[241], tmp18[240], tmp18[239], tmp18[238], tmp18[237], tmp18[236], tmp18[235], tmp18[234], tmp18[233], tmp18[232], tmp18[231], tmp18[230], tmp18[229], tmp18[228], tmp18[227], tmp18[226], tmp18[225], tmp18[224], tmp18[223], tmp18[222], tmp18[221], tmp18[220], tmp18[219], tmp18[218], tmp18[217], tmp18[216], tmp18[215], tmp18[214], tmp18[213], tmp18[212], tmp18[211], tmp18[210], tmp18[209], tmp18[208], tmp18[207], tmp18[206], tmp18[205], tmp18[204], tmp18[203], tmp18[202], tmp18[201], tmp18[200], tmp18[199], tmp18[198], tmp18[197], tmp18[196], tmp18[195], tmp18[194], tmp18[193], tmp18[192], tmp18[191], tmp18[190], tmp18[189], tmp18[188], tmp18[187], tmp18[186], tmp18[185], tmp18[184], tmp18[183], tmp18[182], tmp18[181], tmp18[180], tmp18[179], tmp18[178], tmp18[177], tmp18[176], tmp18[175], tmp18[174], tmp18[173], tmp18[172], tmp18[171], tmp18[170], tmp18[169], tmp18[168], tmp18[167], tmp18[166], tmp18[165], tmp18[164], tmp18[163], tmp18[162], tmp18[161], tmp18[160], tmp18[159], tmp18[158], tmp18[157], tmp18[156], tmp18[155], tmp18[154], tmp18[153], tmp18[152], tmp18[151], tmp18[150], tmp18[149], tmp18[148], tmp18[147], tmp18[146], tmp18[145], tmp18[144], tmp18[143], tmp18[142], tmp18[141], tmp18[140], tmp18[139], tmp18[138], tmp18[137], tmp18[136], tmp18[135], tmp18[134], tmp18[133], tmp18[132], tmp18[131], tmp18[130], tmp18[129], tmp18[128], tmp18[127], tmp18[126], tmp18[125], tmp18[124], tmp18[123], tmp18[122], tmp18[121], tmp18[120], tmp18[119], tmp18[118], tmp18[117], tmp18[116], tmp18[115], tmp18[114], tmp18[113], tmp18[112], tmp18[111], tmp18[110], tmp18[109], tmp18[108], tmp18[107], tmp18[106], tmp18[105], tmp18[104], tmp18[103], tmp18[102], tmp18[101], tmp18[100], tmp18[99], tmp18[98], tmp18[97], tmp18[96], tmp18[95], tmp18[94], tmp18[93], tmp18[92], tmp18[91], tmp18[90], tmp18[89], tmp18[88], tmp18[87], tmp18[86], tmp18[85], tmp18[84], tmp18[83], tmp18[82], tmp18[81], tmp18[80], tmp18[79], tmp18[78], tmp18[77], tmp18[76], tmp18[75], tmp18[74], tmp18[73], tmp18[72], tmp18[71], tmp18[70], tmp18[69], tmp18[68], tmp18[67], tmp18[66], tmp18[65], tmp18[64], tmp18[63], tmp18[62], tmp18[61], tmp18[60], tmp18[59], tmp18[58], tmp18[57], tmp18[56], tmp18[55], tmp18[54], tmp18[53], tmp18[52], tmp18[51], tmp18[50], tmp18[49], tmp18[48], tmp18[47], tmp18[46], tmp18[45], tmp18[44], tmp18[43], tmp18[42], tmp18[41], tmp18[40], tmp18[39], tmp18[38], tmp18[37], tmp18[36], tmp18[35], tmp18[34], tmp18[33], tmp18[32], tmp18[31], tmp18[30], tmp18[29], tmp18[28], tmp18[27], tmp18[26], tmp18[25], tmp18[24], tmp18[23], tmp18[22], tmp18[21], tmp18[20], tmp18[19], tmp18[18], tmp18[17], tmp18[16], tmp18[15], tmp18[14], tmp18[13], tmp18[12], tmp18[11], tmp18[10], tmp18[9], tmp18[8], tmp18[7], tmp18[6], tmp18[5], tmp18[4], tmp18[3], tmp18[2], tmp18[1], tmp18[0]};
    assign tmp7343 = {tmp7342, const_712_0};
    assign tmp7344 = {const_713_0};
    assign tmp7345 = {tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344, tmp7344};
    assign tmp7346 = {tmp7345, const_713_0};
    assign tmp7347 = {tmp18[255]};
    assign tmp7348 = tmp7346 - tmp18;
    assign tmp7349 = {tmp7348[256]};
    assign tmp7350 = {tmp7346[255]};
    assign tmp7351 = ~tmp7350;
    assign tmp7352 = tmp7349 ^ tmp7351;
    assign tmp7353 = {tmp18[255]};
    assign tmp7354 = ~tmp7353;
    assign tmp7355 = tmp7352 ^ tmp7354;
    assign tmp7356 = {tmp7343[255]};
    assign tmp7357 = {const_714_0};
    assign tmp7358 = {tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357, tmp7357};
    assign tmp7359 = {tmp7358, const_714_0};
    assign tmp7360 = tmp7343 - tmp7359;
    assign tmp7361 = {tmp7360[256]};
    assign tmp7362 = {tmp7343[255]};
    assign tmp7363 = ~tmp7362;
    assign tmp7364 = tmp7361 ^ tmp7363;
    assign tmp7365 = {tmp7359[255]};
    assign tmp7366 = ~tmp7365;
    assign tmp7367 = tmp7364 ^ tmp7366;
    assign tmp7368 = tmp7355 & tmp7367;
    assign tmp7369 = {tmp18[255]};
    assign tmp7370 = {const_715_0};
    assign tmp7371 = {tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370, tmp7370};
    assign tmp7372 = {tmp7371, const_715_0};
    assign tmp7373 = tmp18 - tmp7372;
    assign tmp7374 = {tmp7373[256]};
    assign tmp7375 = {tmp18[255]};
    assign tmp7376 = ~tmp7375;
    assign tmp7377 = tmp7374 ^ tmp7376;
    assign tmp7378 = {tmp7372[255]};
    assign tmp7379 = ~tmp7378;
    assign tmp7380 = tmp7377 ^ tmp7379;
    assign tmp7381 = {const_716_0};
    assign tmp7382 = {tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381, tmp7381};
    assign tmp7383 = {tmp7382, const_716_0};
    assign tmp7384 = {tmp7343[255]};
    assign tmp7385 = tmp7383 - tmp7343;
    assign tmp7386 = {tmp7385[256]};
    assign tmp7387 = {tmp7383[255]};
    assign tmp7388 = ~tmp7387;
    assign tmp7389 = tmp7386 ^ tmp7388;
    assign tmp7390 = {tmp7343[255]};
    assign tmp7391 = ~tmp7390;
    assign tmp7392 = tmp7389 ^ tmp7391;
    assign tmp7393 = tmp7383 == tmp7343;
    assign tmp7394 = tmp7392 | tmp7393;
    assign tmp7395 = tmp7380 & tmp7394;
    assign tmp7396 = tmp7368 ? const_717_57896044618658097711785492504343953926634992332820282019728792003956564819967 : tmp7343;
    assign tmp7397 = tmp7395 ? _ver_out_tmp_55 : tmp7396;
    assign tmp7398 = ~tmp35;
    assign tmp7399 = ~tmp36;
    assign tmp7400 = tmp7398 & tmp7399;
    assign tmp7401 = ~tmp57;
    assign tmp7402 = tmp7400 & tmp7401;
    assign tmp7403 = ~tmp1034;
    assign tmp7404 = tmp7402 & tmp7403;
    assign tmp7405 = tmp7404 & tmp2071;
    assign tmp7406 = ~tmp2583;
    assign tmp7407 = tmp7405 & tmp7406;
    assign tmp7408 = ~tmp23;
    assign tmp7409 = tmp7407 & tmp7408;
    assign tmp7410 = tmp7409 & cfg_speculative_egest;
    assign tmp7411 = ~tmp6619;
    assign tmp7412 = tmp7410 & tmp7411;
    assign tmp7413 = tmp7412 & tmp7003;
    assign tmp7414 = ~tmp24;
    assign tmp7415 = tmp7413 & tmp7414;
    assign tmp7416 = ~tmp35;
    assign tmp7417 = ~tmp36;
    assign tmp7418 = tmp7416 & tmp7417;
    assign tmp7419 = ~tmp57;
    assign tmp7420 = tmp7418 & tmp7419;
    assign tmp7421 = ~tmp1034;
    assign tmp7422 = tmp7420 & tmp7421;
    assign tmp7423 = tmp7422 & tmp2071;
    assign tmp7424 = ~tmp2583;
    assign tmp7425 = tmp7423 & tmp7424;
    assign tmp7426 = ~tmp23;
    assign tmp7427 = tmp7425 & tmp7426;
    assign tmp7428 = tmp7427 & cfg_speculative_egest;
    assign tmp7429 = ~tmp6619;
    assign tmp7430 = tmp7428 & tmp7429;
    assign tmp7431 = ~tmp7003;
    assign tmp7432 = tmp7430 & tmp7431;
    assign tmp7433 = ~tmp35;
    assign tmp7434 = ~tmp36;
    assign tmp7435 = tmp7433 & tmp7434;
    assign tmp7436 = ~tmp57;
    assign tmp7437 = tmp7435 & tmp7436;
    assign tmp7438 = ~tmp1034;
    assign tmp7439 = tmp7437 & tmp7438;
    assign tmp7440 = tmp7439 & tmp2071;
    assign tmp7441 = ~tmp2583;
    assign tmp7442 = tmp7440 & tmp7441;
    assign tmp7443 = ~tmp23;
    assign tmp7444 = tmp7442 & tmp7443;
    assign tmp7445 = tmp7444 & cfg_speculative_egest;
    assign tmp7446 = ~tmp6619;
    assign tmp7447 = tmp7445 & tmp7446;
    assign tmp7448 = ~tmp7003;
    assign tmp7449 = tmp7447 & tmp7448;
    assign tmp7450 = ~tmp35;
    assign tmp7451 = ~tmp36;
    assign tmp7452 = tmp7450 & tmp7451;
    assign tmp7453 = ~tmp57;
    assign tmp7454 = tmp7452 & tmp7453;
    assign tmp7455 = ~tmp1034;
    assign tmp7456 = tmp7454 & tmp7455;
    assign tmp7457 = tmp7456 & tmp2071;
    assign tmp7458 = ~tmp2583;
    assign tmp7459 = tmp7457 & tmp7458;
    assign tmp7460 = ~tmp23;
    assign tmp7461 = tmp7459 & tmp7460;
    assign tmp7462 = ~cfg_speculative_egest;
    assign tmp7463 = tmp7461 & tmp7462;
    assign tmp7464 = ~tmp35;
    assign tmp7465 = ~tmp36;
    assign tmp7466 = tmp7464 & tmp7465;
    assign tmp7467 = ~tmp57;
    assign tmp7468 = tmp7466 & tmp7467;
    assign tmp7469 = ~tmp1034;
    assign tmp7470 = tmp7468 & tmp7469;
    assign tmp7471 = tmp7470 & tmp2071;
    assign tmp7472 = ~tmp2583;
    assign tmp7473 = tmp7471 & tmp7472;
    assign tmp7474 = ~tmp23;
    assign tmp7475 = tmp7473 & tmp7474;
    assign tmp7476 = ~cfg_speculative_egest;
    assign tmp7477 = tmp7475 & tmp7476;
    assign tmp7478 = tmp38 ? const_6_0 : tmp11;
    assign tmp7479 = tmp173 ? tmp164 : tmp7478;
    assign tmp7480 = tmp386 ? tmp13 : tmp7479;
    assign tmp7481 = tmp574 ? tmp561 : tmp7480;
    assign tmp7482 = tmp962 ? tmp947 : tmp7481;
    assign tmp7483 = tmp1164 ? tmp1153 : tmp7482;
    assign tmp7484 = tmp1385 ? tmp12 : tmp7483;
    assign tmp7485 = tmp1589 ? tmp1574 : tmp7484;
    assign tmp7486 = tmp1993 ? tmp1976 : tmp7485;
    assign tmp7487 = tmp2671 ? tmp2659 : tmp7486;
    assign tmp7488 = tmp2845 ? tmp2830 : tmp7487;
    assign tmp7489 = tmp2978 ? tmp25 : tmp7488;
    assign tmp7490 = tmp3473 ? tmp29 : tmp7489;
    assign tmp7491 = tmp4074 ? tmp29 : tmp7490;
    assign tmp7492 = tmp4579 ? tmp4557 : tmp7491;
    assign tmp7493 = tmp4768 ? tmp25 : tmp7492;
    assign tmp7494 = tmp5757 ? tmp29 : tmp7493;
    assign tmp7495 = tmp6661 ? tmp15 : tmp7494;
    assign tmp7496 = tmp7056 ? tmp7039 : tmp7495;
    assign tmp7497 = tmp40 ? const_7_2 : tmp12;
    assign tmp7498 = tmp238 ? tmp229 : tmp7497;
    assign tmp7499 = tmp408 ? tmp14 : tmp7498;
    assign tmp7500 = tmp691 ? tmp678 : tmp7499;
    assign tmp7501 = tmp985 ? tmp970 : tmp7500;
    assign tmp7502 = tmp1059 ? tmp11 : tmp7501;
    assign tmp7503 = tmp1398 ? tmp11 : tmp7502;
    assign tmp7504 = tmp1604 ? tmp11 : tmp7503;
    assign tmp7505 = tmp2691 ? tmp2679 : tmp7504;
    assign tmp7506 = tmp2864 ? tmp2849 : tmp7505;
    assign tmp7507 = tmp2994 ? tmp26 : tmp7506;
    assign tmp7508 = tmp3603 ? tmp30 : tmp7507;
    assign tmp7509 = tmp4110 ? tmp30 : tmp7508;
    assign tmp7510 = tmp4605 ? tmp4583 : tmp7509;
    assign tmp7511 = tmp4791 ? tmp26 : tmp7510;
    assign tmp7512 = tmp5901 ? tmp30 : tmp7511;
    assign tmp7513 = tmp6689 ? tmp16 : tmp7512;
    assign tmp7514 = tmp7077 ? tmp7060 : tmp7513;
    assign tmp7515 = tmp42 ? const_8_1 : tmp13;
    assign tmp7516 = tmp76 ? tmp11 : tmp7515;
    assign tmp7517 = tmp397 ? tmp11 : tmp7516;
    assign tmp7518 = tmp587 ? tmp11 : tmp7517;
    assign tmp7519 = tmp1231 ? tmp1220 : tmp7518;
    assign tmp7520 = tmp1411 ? tmp14 : tmp7519;
    assign tmp7521 = tmp1710 ? tmp1695 : tmp7520;
    assign tmp7522 = tmp2018 ? tmp2001 : tmp7521;
    assign tmp7523 = tmp2711 ? tmp2699 : tmp7522;
    assign tmp7524 = tmp2883 ? tmp2868 : tmp7523;
    assign tmp7525 = tmp3010 ? tmp27 : tmp7524;
    assign tmp7526 = tmp3733 ? tmp31 : tmp7525;
    assign tmp7527 = tmp4146 ? tmp31 : tmp7526;
    assign tmp7528 = tmp4631 ? tmp4609 : tmp7527;
    assign tmp7529 = tmp4814 ? tmp27 : tmp7528;
    assign tmp7530 = tmp6045 ? tmp31 : tmp7529;
    assign tmp7531 = tmp6717 ? tmp17 : tmp7530;
    assign tmp7532 = tmp7098 ? tmp7081 : tmp7531;
    assign tmp7533 = tmp44 ? const_9_0 : tmp14;
    assign tmp7534 = tmp83 ? tmp12 : tmp7533;
    assign tmp7535 = tmp419 ? tmp12 : tmp7534;
    assign tmp7536 = tmp704 ? tmp12 : tmp7535;
    assign tmp7537 = tmp1068 ? tmp13 : tmp7536;
    assign tmp7538 = tmp1424 ? tmp13 : tmp7537;
    assign tmp7539 = tmp1725 ? tmp13 : tmp7538;
    assign tmp7540 = tmp2731 ? tmp2719 : tmp7539;
    assign tmp7541 = tmp2902 ? tmp2887 : tmp7540;
    assign tmp7542 = tmp3026 ? tmp28 : tmp7541;
    assign tmp7543 = tmp3863 ? tmp32 : tmp7542;
    assign tmp7544 = tmp4182 ? tmp32 : tmp7543;
    assign tmp7545 = tmp4657 ? tmp4635 : tmp7544;
    assign tmp7546 = tmp4837 ? tmp28 : tmp7545;
    assign tmp7547 = tmp6189 ? tmp32 : tmp7546;
    assign tmp7548 = tmp6745 ? tmp18 : tmp7547;
    assign tmp7549 = tmp7119 ? tmp7102 : tmp7548;
    assign tmp7550 = tmp46 ? const_10_0 : tmp15;
    assign tmp7551 = tmp303 ? tmp294 : tmp7550;
    assign tmp7552 = tmp430 ? tmp17 : tmp7551;
    assign tmp7553 = tmp808 ? tmp795 : tmp7552;
    assign tmp7554 = tmp1008 ? tmp993 : tmp7553;
    assign tmp7555 = tmp1298 ? tmp1287 : tmp7554;
    assign tmp7556 = tmp1437 ? tmp16 : tmp7555;
    assign tmp7557 = tmp1831 ? tmp1816 : tmp7556;
    assign tmp7558 = tmp2043 ? tmp2026 : tmp7557;
    assign tmp7559 = tmp2917 ? tmp29 : tmp7558;
    assign tmp7560 = tmp3098 ? tmp3082 : tmp7559;
    assign tmp7561 = tmp3587 ? tmp3571 : tmp7560;
    assign tmp7562 = tmp4092 ? tmp25 : tmp7561;
    assign tmp7563 = tmp4679 ? tmp29 : tmp7562;
    assign tmp7564 = tmp4916 ? tmp4893 : tmp7563;
    assign tmp7565 = tmp5878 ? tmp5855 : tmp7564;
    assign tmp7566 = tmp6675 ? tmp11 : tmp7565;
    assign tmp7567 = tmp7193 ? tmp7175 : tmp7566;
    assign tmp7568 = tmp48 ? const_11_0 : tmp16;
    assign tmp7569 = tmp368 ? tmp359 : tmp7568;
    assign tmp7570 = tmp452 ? tmp18 : tmp7569;
    assign tmp7571 = tmp925 ? tmp912 : tmp7570;
    assign tmp7572 = tmp1031 ? tmp1016 : tmp7571;
    assign tmp7573 = tmp1077 ? tmp15 : tmp7572;
    assign tmp7574 = tmp1450 ? tmp15 : tmp7573;
    assign tmp7575 = tmp1846 ? tmp15 : tmp7574;
    assign tmp7576 = tmp2932 ? tmp30 : tmp7575;
    assign tmp7577 = tmp3170 ? tmp3154 : tmp7576;
    assign tmp7578 = tmp3717 ? tmp3701 : tmp7577;
    assign tmp7579 = tmp4128 ? tmp26 : tmp7578;
    assign tmp7580 = tmp4701 ? tmp30 : tmp7579;
    assign tmp7581 = tmp4995 ? tmp4972 : tmp7580;
    assign tmp7582 = tmp6022 ? tmp5999 : tmp7581;
    assign tmp7583 = tmp6703 ? tmp12 : tmp7582;
    assign tmp7584 = tmp7267 ? tmp7249 : tmp7583;
    assign tmp7585 = tmp50 ? const_12_0 : tmp17;
    assign tmp7586 = tmp90 ? tmp15 : tmp7585;
    assign tmp7587 = tmp441 ? tmp15 : tmp7586;
    assign tmp7588 = tmp821 ? tmp15 : tmp7587;
    assign tmp7589 = tmp1365 ? tmp1354 : tmp7588;
    assign tmp7590 = tmp1463 ? tmp18 : tmp7589;
    assign tmp7591 = tmp1952 ? tmp1937 : tmp7590;
    assign tmp7592 = tmp2068 ? tmp2051 : tmp7591;
    assign tmp7593 = tmp2947 ? tmp31 : tmp7592;
    assign tmp7594 = tmp3242 ? tmp3226 : tmp7593;
    assign tmp7595 = tmp3847 ? tmp3831 : tmp7594;
    assign tmp7596 = tmp4164 ? tmp27 : tmp7595;
    assign tmp7597 = tmp4723 ? tmp31 : tmp7596;
    assign tmp7598 = tmp5074 ? tmp5051 : tmp7597;
    assign tmp7599 = tmp6166 ? tmp6143 : tmp7598;
    assign tmp7600 = tmp6731 ? tmp13 : tmp7599;
    assign tmp7601 = tmp7341 ? tmp7323 : tmp7600;
    assign tmp7602 = tmp52 ? const_13_1 : tmp18;
    assign tmp7603 = tmp97 ? tmp16 : tmp7602;
    assign tmp7604 = tmp463 ? tmp16 : tmp7603;
    assign tmp7605 = tmp938 ? tmp16 : tmp7604;
    assign tmp7606 = tmp1086 ? tmp17 : tmp7605;
    assign tmp7607 = tmp1476 ? tmp17 : tmp7606;
    assign tmp7608 = tmp1967 ? tmp17 : tmp7607;
    assign tmp7609 = tmp2962 ? tmp32 : tmp7608;
    assign tmp7610 = tmp3314 ? tmp3298 : tmp7609;
    assign tmp7611 = tmp3977 ? tmp3961 : tmp7610;
    assign tmp7612 = tmp4200 ? tmp28 : tmp7611;
    assign tmp7613 = tmp4745 ? tmp32 : tmp7612;
    assign tmp7614 = tmp5153 ? tmp5130 : tmp7613;
    assign tmp7615 = tmp6310 ? tmp6287 : tmp7614;
    assign tmp7616 = tmp6759 ? tmp14 : tmp7615;
    assign tmp7617 = tmp7415 ? tmp7397 : tmp7616;
    assign tmp7618 = tmp54 ? const_14_0 : tmp19;
    assign tmp7619 = tmp65 ? tmp19 : tmp7618;
    assign tmp7620 = tmp1046 ? tmp19 : tmp7619;
    assign tmp7621 = tmp2601 ? const_292_0 : tmp7620;
    assign tmp7622 = tmp2651 ? const_296_0 : tmp7621;
    assign tmp7623 = tmp2826 ? const_318_0 : tmp7622;
    assign tmp7624 = tmp3457 ? const_348_0 : tmp7623;
    assign tmp7625 = tmp4056 ? const_402_0 : tmp7624;
    assign tmp7626 = tmp4553 ? const_432_0 : tmp7625;
    assign tmp7627 = tmp5734 ? const_518_1 : tmp7626;
    assign tmp7628 = tmp6358 ? const_572_0 : tmp7627;
    assign tmp7629 = tmp6400 ? const_574_0 : tmp7628;
    assign tmp7630 = tmp6647 ? const_632_1 : tmp7629;
    assign tmp7631 = tmp7035 ? const_690_1 : tmp7630;
    assign tmp7632 = tmp7449 ? tmp19 : tmp7631;
    assign tmp7633 = tmp7477 ? tmp19 : tmp7632;
    assign tmp7634 = {const_722_0, const_722_0, const_722_0};
    assign tmp7635 = {tmp7634, const_721_0};
    assign tmp7636 = tmp61 ? const_17_0 : tmp7635;
    assign tmp7637 = tmp1040 ? const_118_0 : tmp7636;
    assign tmp7638 = tmp2592 ? const_291_15 : tmp7637;
    assign tmp7639 = tmp2639 ? const_295_8 : tmp7638;
    assign tmp7640 = tmp2812 ? const_317_1 : tmp7639;
    assign tmp7641 = tmp3441 ? const_347_4 : tmp7640;
    assign tmp7642 = tmp4038 ? const_401_6 : tmp7641;
    assign tmp7643 = tmp4532 ? const_431_2 : tmp7642;
    assign tmp7644 = tmp5711 ? const_517_5 : tmp7643;
    assign tmp7645 = tmp6334 ? const_571_0 : tmp7644;
    assign tmp7646 = tmp6379 ? const_573_0 : tmp7645;
    assign tmp7647 = tmp6633 ? const_631_6 : tmp7646;
    assign tmp7648 = tmp7019 ? const_689_3 : tmp7647;
    assign tmp7649 = tmp7432 ? const_719_0 : tmp7648;
    assign tmp7650 = tmp7463 ? const_720_0 : tmp7649;
    assign tmp7651 = tmp2156 ? tmp2148 : const_723_0;
    assign tmp7652 = tmp2241 ? tmp2233 : const_724_0;
    assign tmp7653 = tmp2264 ? tmp2256 : const_725_0;
    assign tmp7654 = tmp2275 ? tmp2267 : const_726_0;
    assign tmp7655 = tmp2291 ? tmp2283 : const_727_0;
    assign tmp7656 = {const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0, const_729_0};
    assign tmp7657 = {tmp7656, const_728_0};
    assign tmp7658 = tmp2334 ? tmp2325 : tmp7657;
    assign tmp7659 = tmp2491 ? tmp11 : tmp7658;
    assign tmp7660 = {const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0, const_731_0};
    assign tmp7661 = {tmp7660, const_730_0};
    assign tmp7662 = tmp2351 ? tmp2342 : tmp7661;
    assign tmp7663 = tmp2502 ? tmp12 : tmp7662;
    assign tmp7664 = {const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0, const_733_0};
    assign tmp7665 = {tmp7664, const_732_0};
    assign tmp7666 = tmp2368 ? tmp2359 : tmp7665;
    assign tmp7667 = tmp2513 ? tmp13 : tmp7666;
    assign tmp7668 = {const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0, const_735_0};
    assign tmp7669 = {tmp7668, const_734_0};
    assign tmp7670 = tmp2385 ? tmp2376 : tmp7669;
    assign tmp7671 = tmp2524 ? tmp14 : tmp7670;
    assign tmp7672 = {const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0, const_737_0};
    assign tmp7673 = {tmp7672, const_736_0};
    assign tmp7674 = tmp2402 ? tmp2393 : tmp7673;
    assign tmp7675 = tmp2535 ? tmp15 : tmp7674;
    assign tmp7676 = {const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0, const_739_0};
    assign tmp7677 = {tmp7676, const_738_0};
    assign tmp7678 = tmp2419 ? tmp2410 : tmp7677;
    assign tmp7679 = tmp2546 ? tmp16 : tmp7678;
    assign tmp7680 = {const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0, const_741_0};
    assign tmp7681 = {tmp7680, const_740_0};
    assign tmp7682 = tmp2436 ? tmp2427 : tmp7681;
    assign tmp7683 = tmp2557 ? tmp17 : tmp7682;
    assign tmp7684 = {const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0, const_743_0};
    assign tmp7685 = {tmp7684, const_742_0};
    assign tmp7686 = tmp2453 ? tmp2444 : tmp7685;
    assign tmp7687 = tmp2568 ? tmp18 : tmp7686;
    assign tmp7689 = {const_745_0, const_745_0};
    assign tmp7690 = {tmp7689, const_744_1};
    assign tmp7691 = tmp7688 == tmp7690;
    assign tmp7692 = {const_747_0};
    assign tmp7693 = {tmp7692, const_746_2};
    assign tmp7694 = tmp7688 == tmp7693;
    assign tmp7695 = tmp7691 | tmp7694;
    assign tmp7696 = {const_749_0};
    assign tmp7697 = {tmp7696, const_748_3};
    assign tmp7698 = tmp7688 == tmp7697;
    assign tmp7699 = tmp7695 | tmp7698;
    assign tmp7700 = {const_751_0};
    assign tmp7701 = {tmp7700, tmp7688};
    assign tmp7702 = tmp7701 == const_750_15;
    assign tmp7703 = tmp7699 | tmp7702;
    assign tmp7704 = tmp7688 == const_752_4;
    assign tmp7705 = tmp7688 == const_753_5;
    assign tmp7706 = tmp7704 | tmp7705;
    assign tmp7707 = tmp7688 == const_754_6;
    assign tmp7708 = tmp7706 | tmp7707;
    assign tmp7709 = tmp7688 == const_755_7;
    assign tmp7710 = tmp7708 | tmp7709;
    assign tmp7711 = {const_757_0};
    assign tmp7712 = {tmp7711, tmp7688};
    assign tmp7713 = tmp7712 == const_756_15;
    assign tmp7714 = tmp7710 | tmp7713;
    assign tmp7715 = {const_759_0};
    assign tmp7716 = {tmp7715, tmp7688};
    assign tmp7717 = tmp7716 == const_758_8;
    assign tmp7718 = tmp7688 == const_760_6;
    assign tmp7719 = tmp7717 | tmp7718;
    assign tmp7720 = tmp7688 == const_761_7;
    assign tmp7721 = tmp7719 | tmp7720;
    assign tmp7722 = {const_763_0};
    assign tmp7723 = {tmp7722, tmp7688};
    assign tmp7724 = tmp7723 == const_762_15;
    assign tmp7725 = tmp7721 | tmp7724;
    assign tmp7726 = {const_765_0, const_765_0};
    assign tmp7727 = {tmp7726, const_764_0};
    assign tmp7728 = my_calculator_ctrl == tmp7727;
    assign tmp7729 = tmp7 & tmp7728;
    assign tmp7730 = {const_768_0, const_768_0};
    assign tmp7731 = {tmp7730, const_767_1};
    assign tmp7732 = my_calculator_ctrl == tmp7731;
    assign tmp7733 = ~tmp7728;
    assign tmp7734 = tmp7 & tmp7733;
    assign tmp7735 = tmp7734 & tmp7732;
    assign tmp7736 = ~tmp7728;
    assign tmp7737 = tmp7 & tmp7736;
    assign tmp7738 = tmp7737 & tmp7732;
    assign tmp7739 = {const_772_0};
    assign tmp7740 = {tmp7739, const_771_2};
    assign tmp7741 = my_calculator_ctrl == tmp7740;
    assign tmp7742 = ~tmp7728;
    assign tmp7743 = tmp7 & tmp7742;
    assign tmp7744 = ~tmp7732;
    assign tmp7745 = tmp7743 & tmp7744;
    assign tmp7746 = tmp7745 & tmp7741;
    assign tmp7747 = ~tmp7728;
    assign tmp7748 = tmp7 & tmp7747;
    assign tmp7749 = ~tmp7732;
    assign tmp7750 = tmp7748 & tmp7749;
    assign tmp7751 = tmp7750 & tmp7741;
    assign tmp7752 = {my_calculator_out_z[2], my_calculator_out_z[1], my_calculator_out_z[0]};
    assign tmp7753 = ~tmp7728;
    assign tmp7754 = tmp7 & tmp7753;
    assign tmp7755 = ~tmp7732;
    assign tmp7756 = tmp7754 & tmp7755;
    assign tmp7757 = tmp7756 & tmp7741;
    assign tmp7758 = {const_776_0};
    assign tmp7759 = {tmp7758, const_775_3};
    assign tmp7760 = my_calculator_ctrl == tmp7759;
    assign tmp7761 = ~tmp7728;
    assign tmp7762 = tmp7 & tmp7761;
    assign tmp7763 = ~tmp7732;
    assign tmp7764 = tmp7762 & tmp7763;
    assign tmp7765 = ~tmp7741;
    assign tmp7766 = tmp7764 & tmp7765;
    assign tmp7767 = tmp7766 & tmp7760;
    assign tmp7768 = {const_779_0, const_779_0};
    assign tmp7769 = {tmp7768, const_778_0};
    assign tmp7770 = tmp7729 ? const_766_1 : tmp7769;
    assign tmp7771 = tmp7738 ? const_770_2 : tmp7770;
    assign tmp7772 = tmp7751 ? const_774_3 : tmp7771;
    assign tmp7773 = tmp7767 ? const_777_1 : tmp7772;
    assign tmp7774 = {const_781_0, const_781_0, const_781_0};
    assign tmp7775 = {tmp7774, const_780_0};
    assign tmp7776 = tmp7735 ? const_769_1 : tmp7775;
    assign tmp7777 = {const_783_0, const_783_0, const_783_0};
    assign tmp7778 = {tmp7777, const_782_0};
    assign tmp7779 = tmp7746 ? const_773_1 : tmp7778;
    assign tmp7780 = tmp7757 ? tmp7752 : tmp7688;

    // Registers
    always @(posedge clk)
    begin
        begin
            tmp0 <= tmp4;
            tmp5 <= tmp6;
            tmp7 <= tmp10;
            tmp11 <= tmp7496;
            tmp12 <= tmp7514;
            tmp13 <= tmp7532;
            tmp14 <= tmp7549;
            tmp15 <= tmp7567;
            tmp16 <= tmp7584;
            tmp17 <= tmp7601;
            tmp18 <= tmp7617;
            tmp19 <= tmp7633;
            tmp7688 <= tmp7780;
        end
    end

endmodule

