// Simple tri-colour LED blink example.

// Correctly map pins for the iCE40UP5K SB_RGBA_DRV hard macro.

`define GREENPWM RGB0PWM
`define REDPWM   RGB1PWM
`define BLUEPWM  RGB2PWM

// taken (mostly) from
// https://github.com/im-tomu/fomu-workshop/blob/master/hdl/verilog/blink-expanded/blink.v

module top (
    // 48MHz Clock input
    // --------
    input clki,
    // LED outputs
    // --------
    output rgb0,
    output rgb1,
    output rgb2,
    // User touchable pins
    // --------
    // Connect 1-2 to enable blue LED
    input  user_1,
    output user_2,
    // Connect 3-4 to enable red LED
    output user_3,
    input  user_4,
    // USB Pins (which should be statically driven if not being used).
    // --------
    output usb_dp,
    output usb_dn,
    output usb_dp_pu
);

    // Assign USB pins to "0" so as to disconnect Fomu from
    // the host system.  Otherwise it would try to talk to
    // us over USB, which wouldn't work since we have no stack.
    assign usb_dp = 1'b0;
    assign usb_dn = 1'b0;
    assign usb_dp_pu = 1'b0;
    // Configure user pins so that we can detect the user connecting
    // 1-2 or 3-4 with conductive material.
    //
    // We do this by grounding user_2 and user_3, and configuring inputs
    // with pullups on user_1 and user_4.
    assign user_2 = 1'b0;
    assign user_3 = 1'b0;

    // Connect to system clock (with buffering)
    wire clk;
    SB_GB clk_gb (
        .USER_SIGNAL_TO_GLOBAL_BUFFER(clki),
        .GLOBAL_BUFFER_OUTPUT(clk)
    );

    // PyRTL module goes here:
    wire [3:0] colors;
    toplevel pyrtl_toplevel (
        .clk (clk),
        .in_1 (~user_1),
        .in_2 (~user_4),
        .red_o (colors[0]),
        .green_o (colors[1]),
        .blue_o (colors[2])
    );

    // Instantiate iCE40 LED driver hard logic, connecting up
    // counter state and LEDs.
    //
    // Note that it's possible to drive the LEDs directly,
    // however that is not current-limited and results in
    // overvolting the red LED.
    //
    // See also:
    // https://www.latticesemi.com/-/media/LatticeSemi/Documents/ApplicationNotes/IK/ICE40LEDDriverUsageGuide.ashx?document_id=50668
    SB_RGBA_DRV #(
        .CURRENT_MODE("0b1"),       // half current
        .RGB0_CURRENT("0b000011"),  // 4 mA
        .RGB1_CURRENT("0b000011"),  // 4 mA
        .RGB2_CURRENT("0b000011")   // 4 mA
    ) RGBA_DRIVER (
        .CURREN(1'b1),
        .RGBLEDEN(1'b1),
        .`REDPWM(colors[0]),      // Red
        .`GREENPWM(colors[1]),    // Green
        .`BLUEPWM(colors[2]),     // Blue
        .RGB0(rgb0),
        .RGB1(rgb1),
        .RGB2(rgb2)
    );

endmodule
// Generated automatically via PyRTL
// As one initial test of synthesis, map to FPGA with:
//   yosys -p "synth_xilinx -top toplevel" thisfile.v

module toplevel(clk, in_1, in_2, blue_o, green_o, red_o);
    input clk;
    input in_1;
    input in_2;
    output blue_o;
    output green_o;
    output red_o;

    reg[2:0] mem_0[31:0]; //tmp7896
    reg[3:0] mem_1[31:0]; //tmp7897
    reg[3:0] mem_2[31:0]; //tmp7898
    reg[2:0] my_calculator_ctrl;
    reg[3:0] my_calculator_in_x;
    reg[3:0] my_calculator_in_y;
    reg[3:0] my_calculator_out_z;
    reg[26:0] tmp0;
    reg tmp5;
    reg tmp7;
    reg[7:0] tmp11;
    reg[7:0] tmp12;
    reg[7:0] tmp13;
    reg[7:0] tmp14;
    reg[7:0] tmp15;
    reg[7:0] tmp16;
    reg[7:0] tmp17;
    reg[7:0] tmp18;
    reg tmp19;
    reg[4:0] tmp7895;
    reg[3:0] tmp7899;

    wire[7:0] _ver_out_tmp_0;
    wire[7:0] _ver_out_tmp_1;
    wire[7:0] _ver_out_tmp_2;
    wire[7:0] _ver_out_tmp_3;
    wire[7:0] _ver_out_tmp_4;
    wire[7:0] _ver_out_tmp_5;
    wire[7:0] _ver_out_tmp_6;
    wire[7:0] _ver_out_tmp_7;
    wire[7:0] _ver_out_tmp_8;
    wire[7:0] _ver_out_tmp_9;
    wire[7:0] _ver_out_tmp_10;
    wire[7:0] _ver_out_tmp_11;
    wire[7:0] _ver_out_tmp_12;
    wire[7:0] _ver_out_tmp_13;
    wire[7:0] _ver_out_tmp_14;
    wire[7:0] _ver_out_tmp_15;
    wire[7:0] _ver_out_tmp_16;
    wire[7:0] _ver_out_tmp_17;
    wire[7:0] _ver_out_tmp_18;
    wire[7:0] _ver_out_tmp_19;
    wire[7:0] _ver_out_tmp_20;
    wire[7:0] _ver_out_tmp_21;
    wire[7:0] _ver_out_tmp_22;
    wire[7:0] _ver_out_tmp_23;
    wire[7:0] _ver_out_tmp_24;
    wire[7:0] _ver_out_tmp_25;
    wire[7:0] _ver_out_tmp_26;
    wire[7:0] _ver_out_tmp_27;
    wire[7:0] _ver_out_tmp_28;
    wire[7:0] _ver_out_tmp_29;
    wire[7:0] _ver_out_tmp_30;
    wire[7:0] _ver_out_tmp_31;
    wire[7:0] _ver_out_tmp_32;
    wire[7:0] _ver_out_tmp_33;
    wire[7:0] _ver_out_tmp_34;
    wire[7:0] _ver_out_tmp_35;
    wire[7:0] _ver_out_tmp_36;
    wire[7:0] _ver_out_tmp_37;
    wire[7:0] _ver_out_tmp_38;
    wire[7:0] _ver_out_tmp_39;
    wire[7:0] _ver_out_tmp_40;
    wire[7:0] _ver_out_tmp_41;
    wire[7:0] _ver_out_tmp_42;
    wire[7:0] _ver_out_tmp_43;
    wire[7:0] _ver_out_tmp_44;
    wire[7:0] _ver_out_tmp_45;
    wire[7:0] _ver_out_tmp_46;
    wire[7:0] _ver_out_tmp_47;
    wire[7:0] _ver_out_tmp_48;
    wire[7:0] _ver_out_tmp_49;
    wire[7:0] _ver_out_tmp_50;
    wire[7:0] _ver_out_tmp_51;
    wire[7:0] _ver_out_tmp_52;
    wire[7:0] _ver_out_tmp_53;
    wire[7:0] _ver_out_tmp_54;
    wire[7:0] _ver_out_tmp_55;
    wire[7:0] _ver_out_tmp_56;
    wire[7:0] _ver_out_tmp_57;
    wire[7:0] _ver_out_tmp_58;
    wire[7:0] _ver_out_tmp_59;
    wire[7:0] _ver_out_tmp_60;
    wire[7:0] _ver_out_tmp_61;
    wire[7:0] _ver_out_tmp_62;
    wire[7:0] _ver_out_tmp_63;
    wire[7:0] _ver_out_tmp_64;
    wire[7:0] _ver_out_tmp_65;
    wire[7:0] _ver_out_tmp_66;
    wire[7:0] _ver_out_tmp_67;
    wire[7:0] _ver_out_tmp_68;
    wire[7:0] _ver_out_tmp_69;
    wire[7:0] _ver_out_tmp_70;
    wire[7:0] _ver_out_tmp_71;
    wire[7:0] _ver_out_tmp_72;
    wire[7:0] _ver_out_tmp_73;
    wire[7:0] _ver_out_tmp_74;
    wire[7:0] _ver_out_tmp_75;
    wire[7:0] _ver_out_tmp_76;
    wire[7:0] _ver_out_tmp_77;
    wire[7:0] _ver_out_tmp_78;
    wire[7:0] _ver_out_tmp_79;
    wire[7:0] _ver_out_tmp_80;
    wire[7:0] _ver_out_tmp_81;
    wire[7:0] _ver_out_tmp_82;
    wire[7:0] _ver_out_tmp_83;
    wire[7:0] _ver_out_tmp_84;
    wire[7:0] _ver_out_tmp_85;
    wire[7:0] _ver_out_tmp_86;
    wire[7:0] _ver_out_tmp_87;
    wire[7:0] _ver_out_tmp_88;
    wire[7:0] _ver_out_tmp_89;
    wire[7:0] _ver_out_tmp_90;
    wire[7:0] _ver_out_tmp_91;
    wire const_1_1;
    wire const_2_0;
    wire const_3_0;
    wire const_4_0;
    wire[2:0] const_5_4;
    wire[7:0] const_6_0;
    wire[7:0] const_7_2;
    wire[7:0] const_8_1;
    wire[7:0] const_9_0;
    wire[7:0] const_10_0;
    wire[7:0] const_11_0;
    wire[7:0] const_12_0;
    wire[7:0] const_13_1;
    wire const_14_0;
    wire const_15_1;
    wire const_16_0;
    wire const_17_0;
    wire const_18_0;
    wire[3:0] const_19_15;
    wire const_20_1;
    wire const_21_0;
    wire[1:0] const_22_2;
    wire const_23_0;
    wire[1:0] const_24_3;
    wire const_25_0;
    wire const_26_0;
    wire const_27_0;
    wire const_28_0;
    wire const_29_0;
    wire const_30_0;
    wire[7:0] const_31_127;
    wire const_33_0;
    wire const_34_0;
    wire const_35_0;
    wire const_36_0;
    wire const_37_0;
    wire[7:0] const_38_127;
    wire const_40_0;
    wire const_41_0;
    wire const_42_0;
    wire const_43_0;
    wire const_44_0;
    wire[7:0] const_45_127;
    wire const_47_0;
    wire const_48_0;
    wire const_49_0;
    wire const_50_0;
    wire const_51_0;
    wire[7:0] const_52_127;
    wire[2:0] const_54_6;
    wire const_55_0;
    wire[2:0] const_56_7;
    wire const_57_0;
    wire[2:0] const_58_4;
    wire const_59_0;
    wire[2:0] const_60_5;
    wire const_61_0;
    wire const_62_0;
    wire const_63_0;
    wire const_64_0;
    wire const_65_0;
    wire const_66_0;
    wire const_67_0;
    wire[7:0] const_68_127;
    wire const_70_0;
    wire const_71_0;
    wire const_72_0;
    wire const_73_0;
    wire const_74_0;
    wire const_75_0;
    wire[7:0] const_76_127;
    wire const_78_0;
    wire const_79_0;
    wire const_80_0;
    wire const_81_0;
    wire const_82_0;
    wire const_83_0;
    wire[7:0] const_84_127;
    wire const_86_0;
    wire const_87_0;
    wire const_88_0;
    wire const_89_0;
    wire const_90_0;
    wire const_91_0;
    wire[7:0] const_92_127;
    wire[3:0] const_94_8;
    wire const_96_0;
    wire const_97_0;
    wire[6:0] const_98_127;
    wire const_99_0;
    wire const_101_0;
    wire const_102_0;
    wire[6:0] const_103_127;
    wire const_104_0;
    wire const_106_0;
    wire const_107_0;
    wire[6:0] const_108_127;
    wire const_109_0;
    wire const_111_0;
    wire const_112_0;
    wire[6:0] const_113_127;
    wire const_114_0;
    wire[1:0] const_115_2;
    wire const_116_0;
    wire const_117_0;
    wire const_118_0;
    wire[3:0] const_119_15;
    wire const_120_1;
    wire const_121_0;
    wire[1:0] const_122_2;
    wire const_123_0;
    wire[1:0] const_124_3;
    wire const_125_0;
    wire const_126_0;
    wire const_127_0;
    wire const_128_0;
    wire const_129_0;
    wire const_130_0;
    wire[7:0] const_131_127;
    wire const_133_0;
    wire const_134_0;
    wire const_135_0;
    wire const_136_0;
    wire const_137_0;
    wire[7:0] const_138_127;
    wire const_140_0;
    wire const_141_0;
    wire const_142_0;
    wire const_143_0;
    wire const_144_0;
    wire[7:0] const_145_127;
    wire const_147_0;
    wire const_148_0;
    wire const_149_0;
    wire const_150_0;
    wire const_151_0;
    wire[7:0] const_152_127;
    wire[2:0] const_154_6;
    wire const_155_0;
    wire[2:0] const_156_7;
    wire const_157_0;
    wire[2:0] const_158_4;
    wire const_159_0;
    wire[2:0] const_160_5;
    wire const_161_0;
    wire const_162_0;
    wire const_163_0;
    wire const_164_0;
    wire const_165_0;
    wire const_166_0;
    wire const_167_0;
    wire[7:0] const_168_127;
    wire const_170_0;
    wire const_171_0;
    wire const_172_0;
    wire const_173_0;
    wire const_174_0;
    wire const_175_0;
    wire[7:0] const_176_127;
    wire const_178_0;
    wire const_179_0;
    wire const_180_0;
    wire const_181_0;
    wire const_182_0;
    wire const_183_0;
    wire[7:0] const_184_127;
    wire const_186_0;
    wire const_187_0;
    wire const_188_0;
    wire const_189_0;
    wire const_190_0;
    wire const_191_0;
    wire[7:0] const_192_127;
    wire[3:0] const_194_8;
    wire const_196_0;
    wire const_197_0;
    wire[6:0] const_198_127;
    wire const_199_0;
    wire const_201_0;
    wire const_202_0;
    wire[6:0] const_203_127;
    wire const_204_0;
    wire const_206_0;
    wire const_207_0;
    wire[6:0] const_208_127;
    wire const_209_0;
    wire const_211_0;
    wire const_212_0;
    wire[6:0] const_213_127;
    wire const_214_0;
    wire[1:0] const_215_3;
    wire const_216_0;
    wire const_217_0;
    wire const_218_0;
    wire const_219_0;
    wire const_220_0;
    wire const_221_0;
    wire const_222_0;
    wire const_223_0;
    wire const_224_0;
    wire const_225_0;
    wire const_226_0;
    wire const_227_0;
    wire const_228_0;
    wire const_229_0;
    wire const_230_0;
    wire const_231_0;
    wire const_232_0;
    wire const_233_0;
    wire const_234_0;
    wire const_235_0;
    wire const_236_0;
    wire const_237_0;
    wire const_238_0;
    wire const_240_0;
    wire const_241_0;
    wire[6:0] const_242_127;
    wire const_243_0;
    wire const_245_0;
    wire const_246_0;
    wire[6:0] const_247_127;
    wire const_248_0;
    wire const_250_0;
    wire const_251_0;
    wire[6:0] const_252_127;
    wire const_253_0;
    wire const_255_0;
    wire const_256_0;
    wire[6:0] const_257_127;
    wire const_258_0;
    wire const_260_0;
    wire const_261_0;
    wire[6:0] const_262_127;
    wire const_263_0;
    wire const_265_0;
    wire const_266_0;
    wire[6:0] const_267_127;
    wire const_268_0;
    wire const_270_0;
    wire const_271_0;
    wire[6:0] const_272_127;
    wire const_273_0;
    wire const_275_0;
    wire const_276_0;
    wire[6:0] const_277_127;
    wire const_278_0;
    wire const_279_0;
    wire const_280_0;
    wire const_281_0;
    wire const_282_0;
    wire const_283_0;
    wire const_284_0;
    wire const_285_0;
    wire const_286_0;
    wire const_287_0;
    wire const_288_0;
    wire[3:0] const_289_15;
    wire const_290_0;
    wire const_291_0;
    wire const_292_0;
    wire[3:0] const_293_8;
    wire const_294_0;
    wire const_296_0;
    wire const_297_0;
    wire[6:0] const_298_127;
    wire const_299_0;
    wire const_301_0;
    wire const_302_0;
    wire[6:0] const_303_127;
    wire const_304_0;
    wire const_306_0;
    wire const_307_0;
    wire[6:0] const_308_127;
    wire const_309_0;
    wire const_311_0;
    wire const_312_0;
    wire[6:0] const_313_127;
    wire const_314_0;
    wire[3:0] const_315_1;
    wire const_316_0;
    wire const_317_0;
    wire const_318_0;
    wire const_319_0;
    wire const_320_0;
    wire const_321_0;
    wire[7:0] const_322_127;
    wire const_324_0;
    wire const_325_0;
    wire const_326_0;
    wire const_327_0;
    wire const_328_0;
    wire[7:0] const_329_127;
    wire const_331_0;
    wire const_332_0;
    wire const_333_0;
    wire const_334_0;
    wire const_335_0;
    wire[7:0] const_336_127;
    wire const_338_0;
    wire const_339_0;
    wire const_340_0;
    wire const_341_0;
    wire const_342_0;
    wire[7:0] const_343_127;
    wire[3:0] const_345_4;
    wire const_346_0;
    wire const_348_0;
    wire const_349_0;
    wire[6:0] const_350_127;
    wire const_351_0;
    wire const_352_0;
    wire const_353_0;
    wire const_354_0;
    wire const_355_0;
    wire const_356_0;
    wire const_357_0;
    wire[7:0] const_358_127;
    wire const_361_0;
    wire const_362_0;
    wire[6:0] const_363_127;
    wire const_364_0;
    wire const_365_0;
    wire const_366_0;
    wire const_367_0;
    wire const_368_0;
    wire const_369_0;
    wire const_370_0;
    wire[7:0] const_371_127;
    wire const_374_0;
    wire const_375_0;
    wire[6:0] const_376_127;
    wire const_377_0;
    wire const_378_0;
    wire const_379_0;
    wire const_380_0;
    wire const_381_0;
    wire const_382_0;
    wire const_383_0;
    wire[7:0] const_384_127;
    wire const_387_0;
    wire const_388_0;
    wire[6:0] const_389_127;
    wire const_390_0;
    wire const_391_0;
    wire const_392_0;
    wire const_393_0;
    wire const_394_0;
    wire const_395_0;
    wire const_396_0;
    wire[7:0] const_397_127;
    wire[3:0] const_399_6;
    wire const_400_0;
    wire[1:0] const_401_0;
    wire const_402_0;
    wire const_403_0;
    wire const_404_0;
    wire const_405_0;
    wire[7:0] const_406_127;
    wire[1:0] const_408_0;
    wire const_409_0;
    wire const_410_0;
    wire const_411_0;
    wire const_412_0;
    wire[7:0] const_413_127;
    wire[1:0] const_415_0;
    wire const_416_0;
    wire const_417_0;
    wire const_418_0;
    wire const_419_0;
    wire[7:0] const_420_127;
    wire[1:0] const_422_0;
    wire const_423_0;
    wire const_424_0;
    wire const_425_0;
    wire const_426_0;
    wire[7:0] const_427_127;
    wire[3:0] const_429_2;
    wire const_430_0;
    wire const_431_0;
    wire const_432_0;
    wire const_433_0;
    wire const_434_0;
    wire const_435_0;
    wire[7:0] const_436_127;
    wire const_438_0;
    wire const_439_0;
    wire const_440_0;
    wire const_441_0;
    wire const_442_0;
    wire[7:0] const_443_127;
    wire const_445_0;
    wire const_446_0;
    wire const_447_0;
    wire const_448_0;
    wire const_449_0;
    wire[7:0] const_450_127;
    wire const_452_0;
    wire const_453_0;
    wire const_454_0;
    wire const_455_0;
    wire const_456_0;
    wire[7:0] const_457_127;
    wire const_459_0;
    wire const_460_0;
    wire const_461_0;
    wire const_462_0;
    wire const_463_0;
    wire[7:0] const_464_127;
    wire const_466_0;
    wire const_467_0;
    wire const_468_0;
    wire const_469_0;
    wire const_470_0;
    wire[7:0] const_471_127;
    wire const_473_0;
    wire const_474_0;
    wire const_475_0;
    wire const_476_0;
    wire const_477_0;
    wire[7:0] const_478_127;
    wire const_480_0;
    wire const_481_0;
    wire const_482_0;
    wire const_483_0;
    wire const_484_0;
    wire[7:0] const_485_127;
    wire const_487_0;
    wire const_488_0;
    wire const_489_0;
    wire const_490_0;
    wire const_491_0;
    wire[7:0] const_492_127;
    wire const_494_0;
    wire const_495_0;
    wire const_496_0;
    wire const_497_0;
    wire const_498_0;
    wire[7:0] const_499_127;
    wire const_501_0;
    wire const_502_0;
    wire const_503_0;
    wire const_504_0;
    wire const_505_0;
    wire[7:0] const_506_127;
    wire const_508_0;
    wire const_509_0;
    wire const_510_0;
    wire const_511_0;
    wire const_512_0;
    wire[7:0] const_513_127;
    wire[3:0] const_515_5;
    wire const_516_1;
    wire const_518_0;
    wire const_519_0;
    wire[6:0] const_520_127;
    wire const_521_0;
    wire const_522_0;
    wire const_523_0;
    wire const_524_0;
    wire const_525_0;
    wire const_526_0;
    wire const_527_0;
    wire[7:0] const_528_127;
    wire const_531_0;
    wire const_532_0;
    wire[6:0] const_533_127;
    wire const_534_0;
    wire const_535_0;
    wire const_536_0;
    wire const_537_0;
    wire const_538_0;
    wire const_539_0;
    wire const_540_0;
    wire[7:0] const_541_127;
    wire const_544_0;
    wire const_545_0;
    wire[6:0] const_546_127;
    wire const_547_0;
    wire const_548_0;
    wire const_549_0;
    wire const_550_0;
    wire const_551_0;
    wire const_552_0;
    wire const_553_0;
    wire[7:0] const_554_127;
    wire const_557_0;
    wire const_558_0;
    wire[6:0] const_559_127;
    wire const_560_0;
    wire const_561_0;
    wire const_562_0;
    wire const_563_0;
    wire const_564_0;
    wire const_565_0;
    wire const_566_0;
    wire[7:0] const_567_127;
    wire[3:0] const_569_0;
    wire const_570_0;
    wire[3:0] const_571_0;
    wire const_572_0;
    wire const_573_1;
    wire const_575_0;
    wire const_576_0;
    wire[6:0] const_577_127;
    wire const_578_0;
    wire const_579_0;
    wire const_580_1;
    wire const_582_0;
    wire const_583_0;
    wire[6:0] const_584_127;
    wire const_585_0;
    wire const_586_0;
    wire const_587_1;
    wire const_589_0;
    wire const_590_0;
    wire[6:0] const_591_127;
    wire const_592_0;
    wire const_593_0;
    wire const_594_1;
    wire const_596_0;
    wire const_597_0;
    wire[6:0] const_598_127;
    wire const_599_0;
    wire const_600_0;
    wire const_601_1;
    wire const_603_0;
    wire const_604_0;
    wire[6:0] const_605_127;
    wire const_606_0;
    wire const_607_0;
    wire const_608_1;
    wire const_610_0;
    wire const_611_0;
    wire[6:0] const_612_127;
    wire const_613_0;
    wire const_614_0;
    wire const_615_1;
    wire const_617_0;
    wire const_618_0;
    wire[6:0] const_619_127;
    wire const_620_0;
    wire const_621_0;
    wire const_622_1;
    wire const_624_0;
    wire const_625_0;
    wire[6:0] const_626_127;
    wire const_627_0;
    wire const_628_0;
    wire[3:0] const_629_7;
    wire const_630_1;
    wire const_631_1;
    wire const_633_0;
    wire const_634_0;
    wire[6:0] const_635_127;
    wire const_636_0;
    wire const_637_0;
    wire const_638_1;
    wire const_640_0;
    wire const_641_0;
    wire[6:0] const_642_127;
    wire const_643_0;
    wire const_644_0;
    wire const_645_1;
    wire const_647_0;
    wire const_648_0;
    wire[6:0] const_649_127;
    wire const_650_0;
    wire const_651_0;
    wire const_652_1;
    wire const_654_0;
    wire const_655_0;
    wire[6:0] const_656_127;
    wire const_657_0;
    wire const_658_0;
    wire const_659_1;
    wire const_661_0;
    wire const_662_0;
    wire[6:0] const_663_127;
    wire const_664_0;
    wire const_665_0;
    wire const_666_1;
    wire const_668_0;
    wire const_669_0;
    wire[6:0] const_670_127;
    wire const_671_0;
    wire const_672_0;
    wire const_673_1;
    wire const_675_0;
    wire const_676_0;
    wire[6:0] const_677_127;
    wire const_678_0;
    wire const_679_0;
    wire const_680_1;
    wire const_682_0;
    wire const_683_0;
    wire[6:0] const_684_127;
    wire const_685_0;
    wire const_686_0;
    wire[3:0] const_687_3;
    wire const_688_1;
    wire const_689_0;
    wire const_690_0;
    wire const_691_0;
    wire const_692_0;
    wire const_693_0;
    wire[7:0] const_694_127;
    wire const_696_0;
    wire const_697_0;
    wire const_698_0;
    wire const_699_0;
    wire const_700_0;
    wire[7:0] const_701_127;
    wire const_703_0;
    wire const_704_0;
    wire const_705_0;
    wire const_706_0;
    wire const_707_0;
    wire[7:0] const_708_127;
    wire const_710_0;
    wire const_711_0;
    wire const_712_0;
    wire const_713_0;
    wire const_714_0;
    wire[7:0] const_715_127;
    wire[3:0] const_717_0;
    wire[3:0] const_718_0;
    wire const_719_0;
    wire const_720_0;
    wire const_721_0;
    wire const_722_0;
    wire const_723_0;
    wire const_724_0;
    wire const_725_0;
    wire const_726_0;
    wire const_727_0;
    wire const_728_0;
    wire const_729_0;
    wire const_730_0;
    wire const_731_0;
    wire const_732_0;
    wire const_733_0;
    wire const_734_0;
    wire const_735_0;
    wire const_736_0;
    wire const_737_0;
    wire const_738_0;
    wire const_739_0;
    wire const_740_1;
    wire const_741_0;
    wire[1:0] const_742_2;
    wire const_743_0;
    wire[1:0] const_744_3;
    wire const_745_0;
    wire[3:0] const_746_15;
    wire[2:0] const_747_4;
    wire const_748_0;
    wire[2:0] const_749_5;
    wire const_750_0;
    wire[2:0] const_751_6;
    wire const_752_0;
    wire[2:0] const_753_7;
    wire const_754_0;
    wire[3:0] const_755_15;
    wire[3:0] const_756_8;
    wire[2:0] const_757_6;
    wire const_758_0;
    wire[2:0] const_759_7;
    wire const_760_0;
    wire[3:0] const_761_15;
    wire const_762_1;
    wire const_763_0;
    wire[2:0] const_764_4;
    wire[3:0] const_765_8;
    wire const_766_1;
    wire const_767_0;
    wire[1:0] const_768_2;
    wire const_769_0;
    wire[3:0] const_770_6;
    wire[1:0] const_771_3;
    wire const_772_0;
    wire[3:0] const_773_6;
    wire const_778_0;
    wire const_779_0;
    wire const_780_0;
    wire const_781_0;
    wire[25:0] tmp1;
    wire[26:0] tmp2;
    wire[27:0] tmp3;
    wire[26:0] tmp4;
    wire tmp8;
    wire tmp9;
    wire tmp10;
    wire tmp33;
    wire[2:0] tmp35;
    wire tmp36;
    wire tmp37;
    wire tmp61;
    wire[2:0] tmp75;
    wire tmp76;
    wire tmp85;
    wire tmp86;
    wire tmp94;
    wire tmp122;
    wire tmp125;
    wire tmp128;
    wire tmp129;
    wire tmp132;
    wire tmp133;
    wire tmp146;
    wire tmp156;
    wire tmp160;
    wire tmp171;
    wire[8:0] tmp177;
    wire tmp178;
    wire tmp186;
    wire tmp187;
    wire tmp196;
    wire[6:0] tmp201;
    wire[7:0] tmp202;
    wire tmp214;
    wire[8:0] tmp219;
    wire tmp220;
    wire tmp222;
    wire tmp223;
    wire tmp226;
    wire tmp227;
    wire[8:0] tmp232;
    wire tmp235;
    wire[8:0] tmp244;
    wire tmp245;
    wire tmp248;
    wire tmp249;
    wire tmp251;
    wire tmp252;
    wire tmp253;
    wire tmp254;
    wire[7:0] tmp255;
    wire[7:0] tmp256;
    wire[6:0] tmp268;
    wire tmp287;
    wire tmp290;
    wire[8:0] tmp299;
    wire tmp312;
    wire tmp320;
    wire tmp334;
    wire tmp345;
    wire tmp354;
    wire tmp388;
    wire tmp404;
    wire tmp407;
    wire tmp408;
    wire tmp421;
    wire tmp444;
    wire tmp445;
    wire[3:0] tmp514;
    wire tmp515;
    wire tmp518;
    wire tmp519;
    wire tmp520;
    wire[9:0] tmp526;
    wire[8:0] tmp527;
    wire[7:0] tmp528;
    wire tmp549;
    wire tmp550;
    wire tmp553;
    wire[8:0] tmp558;
    wire tmp559;
    wire tmp562;
    wire tmp565;
    wire tmp566;
    wire tmp567;
    wire tmp568;
    wire[8:0] tmp573;
    wire tmp592;
    wire tmp593;
    wire[8:0] tmp598;
    wire tmp599;
    wire tmp602;
    wire tmp603;
    wire tmp604;
    wire tmp605;
    wire tmp607;
    wire tmp608;
    wire[7:0] tmp609;
    wire[7:0] tmp610;
    wire tmp644;
    wire[8:0] tmp646;
    wire[9:0] tmp647;
    wire[8:0] tmp648;
    wire[7:0] tmp649;
    wire tmp674;
    wire[8:0] tmp679;
    wire tmp680;
    wire tmp681;
    wire tmp682;
    wire tmp683;
    wire tmp686;
    wire tmp687;
    wire tmp688;
    wire tmp689;
    wire tmp698;
    wire tmp701;
    wire tmp714;
    wire[8:0] tmp719;
    wire tmp720;
    wire tmp723;
    wire tmp726;
    wire tmp728;
    wire tmp729;
    wire[7:0] tmp730;
    wire[7:0] tmp731;
    wire[9:0] tmp768;
    wire[8:0] tmp769;
    wire[7:0] tmp770;
    wire tmp795;
    wire[8:0] tmp800;
    wire tmp801;
    wire tmp803;
    wire tmp804;
    wire tmp807;
    wire tmp808;
    wire tmp809;
    wire tmp810;
    wire tmp819;
    wire tmp835;
    wire[8:0] tmp840;
    wire tmp841;
    wire tmp844;
    wire tmp845;
    wire tmp847;
    wire tmp849;
    wire tmp850;
    wire[7:0] tmp851;
    wire[7:0] tmp852;
    wire[8:0] tmp888;
    wire[9:0] tmp889;
    wire[8:0] tmp890;
    wire[7:0] tmp891;
    wire tmp897;
    wire tmp902;
    wire tmp909;
    wire tmp912;
    wire tmp916;
    wire[8:0] tmp921;
    wire tmp922;
    wire tmp923;
    wire tmp924;
    wire tmp925;
    wire tmp928;
    wire tmp930;
    wire tmp931;
    wire tmp937;
    wire tmp938;
    wire tmp956;
    wire[8:0] tmp961;
    wire tmp962;
    wire tmp965;
    wire tmp968;
    wire tmp969;
    wire tmp970;
    wire tmp971;
    wire[7:0] tmp972;
    wire[7:0] tmp973;
    wire tmp988;
    wire tmp1004;
    wire tmp1005;
    wire tmp1028;
    wire tmp1030;
    wire tmp1046;
    wire[7:0] tmp1062;
    wire tmp1077;
    wire tmp1093;
    wire tmp1099;
    wire tmp1100;
    wire tmp1101;
    wire tmp1104;
    wire[2:0] tmp1106;
    wire tmp1107;
    wire tmp1111;
    wire[3:0] tmp1117;
    wire tmp1118;
    wire tmp1119;
    wire tmp1127;
    wire tmp1141;
    wire[2:0] tmp1164;
    wire[3:0] tmp1165;
    wire tmp1166;
    wire tmp1169;
    wire tmp1170;
    wire tmp1173;
    wire tmp1174;
    wire[6:0] tmp1175;
    wire[7:0] tmp1176;
    wire[8:0] tmp1181;
    wire tmp1182;
    wire[8:0] tmp1193;
    wire tmp1194;
    wire tmp1196;
    wire tmp1200;
    wire tmp1222;
    wire tmp1223;
    wire tmp1225;
    wire tmp1226;
    wire[7:0] tmp1229;
    wire[7:0] tmp1230;
    wire tmp1240;
    wire[6:0] tmp1244;
    wire[7:0] tmp1245;
    wire[8:0] tmp1250;
    wire tmp1251;
    wire[8:0] tmp1262;
    wire tmp1263;
    wire tmp1264;
    wire tmp1266;
    wire tmp1269;
    wire tmp1270;
    wire tmp1279;
    wire[8:0] tmp1287;
    wire tmp1288;
    wire tmp1291;
    wire tmp1293;
    wire tmp1294;
    wire tmp1295;
    wire tmp1296;
    wire tmp1297;
    wire[7:0] tmp1298;
    wire[7:0] tmp1299;
    wire tmp1320;
    wire tmp1326;
    wire[8:0] tmp1331;
    wire tmp1338;
    wire tmp1361;
    wire tmp1362;
    wire tmp1363;
    wire[7:0] tmp1367;
    wire tmp1381;
    wire tmp1392;
    wire[8:0] tmp1400;
    wire tmp1404;
    wire tmp1407;
    wire[8:0] tmp1413;
    wire tmp1420;
    wire[8:0] tmp1425;
    wire tmp1426;
    wire tmp1429;
    wire tmp1434;
    wire tmp1435;
    wire[7:0] tmp1436;
    wire[7:0] tmp1437;
    wire[3:0] tmp1452;
    wire tmp1453;
    wire[3:0] tmp1455;
    wire tmp1456;
    wire tmp1457;
    wire tmp1468;
    wire tmp1496;
    wire tmp1548;
    wire tmp1577;
    wire tmp1580;
    wire tmp1583;
    wire tmp1584;
    wire[8:0] tmp1587;
    wire[8:0] tmp1590;
    wire[9:0] tmp1591;
    wire[8:0] tmp1592;
    wire[7:0] tmp1593;
    wire tmp1602;
    wire tmp1605;
    wire tmp1611;
    wire tmp1614;
    wire tmp1615;
    wire tmp1618;
    wire[8:0] tmp1623;
    wire tmp1624;
    wire tmp1625;
    wire tmp1626;
    wire tmp1627;
    wire tmp1630;
    wire tmp1632;
    wire tmp1633;
    wire tmp1658;
    wire[8:0] tmp1663;
    wire tmp1664;
    wire tmp1667;
    wire tmp1670;
    wire tmp1671;
    wire tmp1672;
    wire tmp1673;
    wire[7:0] tmp1674;
    wire[7:0] tmp1675;
    wire tmp1709;
    wire[8:0] tmp1712;
    wire[9:0] tmp1716;
    wire[8:0] tmp1717;
    wire[7:0] tmp1718;
    wire tmp1730;
    wire[8:0] tmp1735;
    wire tmp1736;
    wire tmp1739;
    wire tmp1742;
    wire tmp1743;
    wire[8:0] tmp1748;
    wire tmp1749;
    wire tmp1750;
    wire tmp1752;
    wire tmp1755;
    wire tmp1756;
    wire tmp1757;
    wire tmp1758;
    wire[8:0] tmp1763;
    wire tmp1764;
    wire tmp1776;
    wire tmp1778;
    wire tmp1783;
    wire[8:0] tmp1788;
    wire tmp1789;
    wire tmp1792;
    wire tmp1794;
    wire tmp1795;
    wire tmp1797;
    wire tmp1798;
    wire[7:0] tmp1799;
    wire[7:0] tmp1800;
    wire tmp1815;
    wire[8:0] tmp1837;
    wire[8:0] tmp1840;
    wire[9:0] tmp1841;
    wire[8:0] tmp1842;
    wire[7:0] tmp1843;
    wire[8:0] tmp1860;
    wire tmp1868;
    wire[8:0] tmp1873;
    wire tmp1874;
    wire tmp1876;
    wire tmp1877;
    wire tmp1880;
    wire tmp1882;
    wire tmp1883;
    wire tmp1889;
    wire tmp1904;
    wire tmp1908;
    wire[8:0] tmp1913;
    wire tmp1914;
    wire tmp1917;
    wire tmp1918;
    wire tmp1920;
    wire tmp1921;
    wire tmp1922;
    wire tmp1923;
    wire[7:0] tmp1924;
    wire[7:0] tmp1925;
    wire[8:0] tmp1962;
    wire[9:0] tmp1966;
    wire[8:0] tmp1967;
    wire[7:0] tmp1968;
    wire[8:0] tmp1973;
    wire tmp1979;
    wire tmp1980;
    wire tmp1993;
    wire[8:0] tmp1998;
    wire tmp1999;
    wire tmp2000;
    wire tmp2001;
    wire tmp2002;
    wire tmp2005;
    wire tmp2007;
    wire tmp2008;
    wire tmp2014;
    wire tmp2026;
    wire tmp2032;
    wire tmp2033;
    wire[8:0] tmp2038;
    wire tmp2039;
    wire tmp2042;
    wire tmp2045;
    wire tmp2046;
    wire tmp2047;
    wire tmp2048;
    wire[7:0] tmp2049;
    wire[7:0] tmp2050;
    wire tmp2085;
    wire tmp2095;
    wire tmp2113;
    wire[7:0] tmp2120;
    wire tmp2138;
    wire tmp2159;
    wire tmp2164;
    wire[7:0] tmp2174;
    wire tmp2187;
    wire tmp2188;
    wire tmp2190;
    wire tmp2193;
    wire[2:0] tmp2195;
    wire tmp2196;
    wire tmp2214;
    wire tmp2221;
    wire tmp2246;
    wire tmp2247;
    wire tmp2255;
    wire[8:0] tmp2264;
    wire tmp2268;
    wire tmp2271;
    wire tmp2272;
    wire tmp2273;
    wire tmp2308;
    wire tmp2320;
    wire tmp2333;
    wire tmp2334;
    wire[8:0] tmp2351;
    wire tmp2354;
    wire tmp2355;
    wire tmp2359;
    wire tmp2360;
    wire tmp2377;
    wire tmp2380;
    wire tmp2381;
    wire tmp2384;
    wire tmp2385;
    wire tmp2396;
    wire tmp2397;
    wire tmp2398;
    wire tmp2409;
    wire tmp2410;
    wire tmp2411;
    wire tmp2412;
    wire tmp2413;
    wire tmp2414;
    wire tmp2415;
    wire tmp2416;
    wire tmp2432;
    wire tmp2439;
    wire tmp2452;
    wire[8:0] tmp2459;
    wire[7:0] tmp2460;
    wire[8:0] tmp2516;
    wire[7:0] tmp2517;
    wire[8:0] tmp2534;
    wire tmp2548;
    wire[7:0] tmp2555;
    wire tmp2566;
    wire tmp2586;
    wire[7:0] tmp2593;
    wire tmp2623;
    wire tmp2628;
    wire tmp2629;
    wire tmp2630;
    wire tmp2631;
    wire tmp2702;
    wire tmp2706;
    wire tmp2730;
    wire tmp2733;
    wire tmp2734;
    wire tmp2735;
    wire[6:0] tmp2736;
    wire tmp2738;
    wire tmp2741;
    wire tmp2742;
    wire tmp2746;
    wire tmp2750;
    wire tmp2772;
    wire tmp2781;
    wire tmp2784;
    wire tmp2797;
    wire tmp2798;
    wire[7:0] tmp2856;
    wire[8:0] tmp2877;
    wire tmp2892;
    wire tmp2916;
    wire[8:0] tmp2921;
    wire tmp2922;
    wire tmp2923;
    wire tmp2924;
    wire tmp2925;
    wire tmp2928;
    wire tmp2929;
    wire tmp2930;
    wire[8:0] tmp2937;
    wire tmp2938;
    wire tmp2941;
    wire tmp2944;
    wire tmp2945;
    wire tmp2946;
    wire tmp2947;
    wire[6:0] tmp2948;
    wire[8:0] tmp2954;
    wire tmp2955;
    wire tmp2958;
    wire tmp2961;
    wire tmp2962;
    wire tmp2963;
    wire tmp2964;
    wire[8:0] tmp2971;
    wire tmp2972;
    wire tmp2974;
    wire tmp2975;
    wire tmp2978;
    wire tmp2979;
    wire tmp2980;
    wire tmp2981;
    wire tmp3036;
    wire[7:0] tmp3038;
    wire tmp3055;
    wire[6:0] tmp3077;
    wire tmp3078;
    wire tmp3113;
    wire tmp3157;
    wire tmp3194;
    wire tmp3197;
    wire tmp3201;
    wire[6:0] tmp3238;
    wire[7:0] tmp3239;
    wire tmp3245;
    wire tmp3260;
    wire tmp3270;
    wire tmp3282;
    wire tmp3285;
    wire tmp3286;
    wire tmp3288;
    wire tmp3290;
    wire tmp3291;
    wire tmp3298;
    wire tmp3319;
    wire tmp3322;
    wire tmp3350;
    wire[7:0] tmp3366;
    wire[7:0] tmp3367;
    wire[8:0] tmp3404;
    wire[8:0] tmp3417;
    wire tmp3421;
    wire[8:0] tmp3429;
    wire tmp3430;
    wire tmp3433;
    wire tmp3435;
    wire tmp3436;
    wire tmp3438;
    wire[7:0] tmp3440;
    wire[6:0] tmp3460;
    wire[7:0] tmp3461;
    wire tmp3470;
    wire tmp3473;
    wire tmp3486;
    wire[8:0] tmp3491;
    wire tmp3492;
    wire tmp3495;
    wire tmp3498;
    wire tmp3504;
    wire tmp3507;
    wire tmp3511;
    wire tmp3512;
    wire[7:0] tmp3515;
    wire tmp3537;
    wire tmp3540;
    wire tmp3543;
    wire tmp3544;
    wire tmp3545;
    wire tmp3551;
    wire tmp3552;
    wire tmp3554;
    wire tmp3555;
    wire tmp3556;
    wire tmp3557;
    wire tmp3558;
    wire tmp3562;
    wire tmp3565;
    wire tmp3568;
    wire tmp3569;
    wire tmp3570;
    wire tmp3571;
    wire[8:0] tmp3574;
    wire tmp3575;
    wire tmp3578;
    wire tmp3579;
    wire tmp3581;
    wire tmp3582;
    wire tmp3583;
    wire tmp3584;
    wire[7:0] tmp3588;
    wire[8:0] tmp3591;
    wire tmp3592;
    wire tmp3595;
    wire tmp3598;
    wire tmp3599;
    wire[8:0] tmp3606;
    wire tmp3607;
    wire tmp3608;
    wire tmp3609;
    wire tmp3610;
    wire tmp3613;
    wire tmp3614;
    wire[8:0] tmp3621;
    wire tmp3622;
    wire tmp3623;
    wire tmp3624;
    wire tmp3625;
    wire tmp3628;
    wire tmp3629;
    wire[7:0] tmp3633;
    wire[8:0] tmp3636;
    wire tmp3637;
    wire tmp3638;
    wire tmp3640;
    wire tmp3643;
    wire tmp3644;
    wire tmp3698;
    wire tmp3699;
    wire[8:0] tmp3705;
    wire[9:0] tmp3708;
    wire[9:0] tmp3711;
    wire[10:0] tmp3712;
    wire[9:0] tmp3713;
    wire[9:0] tmp3731;
    wire tmp3732;
    wire tmp3735;
    wire tmp3736;
    wire tmp3737;
    wire tmp3738;
    wire tmp3739;
    wire tmp3746;
    wire tmp3747;
    wire tmp3748;
    wire tmp3752;
    wire tmp3753;
    wire tmp3754;
    wire[8:0] tmp3759;
    wire tmp3760;
    wire tmp3762;
    wire[9:0] tmp3771;
    wire tmp3775;
    wire tmp3794;
    wire[7:0] tmp3795;
    wire tmp3833;
    wire[1:0] tmp3841;
    wire[9:0] tmp3842;
    wire[9:0] tmp3845;
    wire[10:0] tmp3846;
    wire[8:0] tmp3853;
    wire tmp3854;
    wire tmp3857;
    wire[9:0] tmp3865;
    wire[8:0] tmp3878;
    wire[8:0] tmp3893;
    wire tmp3894;
    wire tmp3895;
    wire tmp3897;
    wire tmp3906;
    wire tmp3925;
    wire tmp3927;
    wire tmp3928;
    wire[8:0] tmp3970;
    wire[8:0] tmp3973;
    wire[1:0] tmp3975;
    wire[9:0] tmp3976;
    wire[9:0] tmp3979;
    wire tmp3994;
    wire[9:0] tmp3999;
    wire tmp4003;
    wire tmp4005;
    wire tmp4007;
    wire tmp4021;
    wire tmp4040;
    wire tmp4041;
    wire tmp4043;
    wire tmp4046;
    wire tmp4047;
    wire tmp4053;
    wire tmp4060;
    wire[7:0] tmp4064;
    wire tmp4101;
    wire[9:0] tmp4113;
    wire[7:0] tmp4116;
    wire[8:0] tmp4121;
    wire tmp4122;
    wire tmp4125;
    wire tmp4134;
    wire[8:0] tmp4146;
    wire tmp4147;
    wire tmp4149;
    wire tmp4163;
    wire tmp4164;
    wire tmp4174;
    wire tmp4180;
    wire tmp4187;
    wire tmp4191;
    wire tmp4194;
    wire[7:0] tmp4198;
    wire[8:0] tmp4219;
    wire tmp4220;
    wire tmp4223;
    wire tmp4226;
    wire[8:0] tmp4229;
    wire tmp4230;
    wire tmp4233;
    wire tmp4236;
    wire tmp4237;
    wire[8:0] tmp4240;
    wire tmp4241;
    wire tmp4244;
    wire tmp4246;
    wire tmp4247;
    wire tmp4248;
    wire[8:0] tmp4251;
    wire tmp4252;
    wire tmp4255;
    wire tmp4258;
    wire tmp4259;
    wire tmp4274;
    wire tmp4311;
    wire tmp4359;
    wire tmp4442;
    wire tmp4456;
    wire[8:0] tmp4462;
    wire tmp4466;
    wire tmp4469;
    wire[5:0] tmp4470;
    wire[7:0] tmp4471;
    wire[8:0] tmp4488;
    wire tmp4489;
    wire tmp4490;
    wire tmp4492;
    wire tmp4495;
    wire tmp4496;
    wire[8:0] tmp4513;
    wire tmp4514;
    wire tmp4517;
    wire tmp4519;
    wire tmp4520;
    wire tmp4521;
    wire tmp4522;
    wire tmp4523;
    wire[7:0] tmp4524;
    wire[7:0] tmp4525;
    wire[8:0] tmp4528;
    wire tmp4529;
    wire tmp4532;
    wire tmp4533;
    wire tmp4534;
    wire tmp4535;
    wire tmp4536;
    wire[8:0] tmp4539;
    wire tmp4540;
    wire tmp4543;
    wire tmp4546;
    wire tmp4547;
    wire[5:0] tmp4548;
    wire[7:0] tmp4549;
    wire tmp4561;
    wire[8:0] tmp4566;
    wire tmp4567;
    wire tmp4568;
    wire tmp4569;
    wire tmp4570;
    wire tmp4573;
    wire tmp4574;
    wire tmp4583;
    wire[8:0] tmp4591;
    wire tmp4592;
    wire tmp4595;
    wire tmp4598;
    wire tmp4599;
    wire tmp4600;
    wire tmp4601;
    wire[7:0] tmp4602;
    wire[7:0] tmp4603;
    wire[8:0] tmp4606;
    wire tmp4607;
    wire tmp4610;
    wire tmp4611;
    wire tmp4612;
    wire tmp4613;
    wire tmp4614;
    wire[8:0] tmp4617;
    wire tmp4619;
    wire tmp4621;
    wire tmp4623;
    wire tmp4624;
    wire tmp4625;
    wire[5:0] tmp4626;
    wire[7:0] tmp4627;
    wire tmp4633;
    wire[8:0] tmp4644;
    wire tmp4645;
    wire tmp4646;
    wire tmp4648;
    wire tmp4651;
    wire tmp4652;
    wire[8:0] tmp4669;
    wire tmp4670;
    wire tmp4673;
    wire tmp4675;
    wire tmp4676;
    wire tmp4677;
    wire tmp4678;
    wire tmp4679;
    wire[7:0] tmp4680;
    wire[7:0] tmp4681;
    wire[8:0] tmp4684;
    wire tmp4685;
    wire tmp4688;
    wire tmp4689;
    wire tmp4690;
    wire tmp4691;
    wire tmp4692;
    wire tmp4698;
    wire tmp4699;
    wire tmp4702;
    wire tmp4703;
    wire[5:0] tmp4704;
    wire[7:0] tmp4705;
    wire tmp4711;
    wire[8:0] tmp4722;
    wire tmp4723;
    wire tmp4724;
    wire tmp4725;
    wire tmp4726;
    wire tmp4729;
    wire tmp4730;
    wire[8:0] tmp4747;
    wire tmp4748;
    wire tmp4751;
    wire tmp4754;
    wire tmp4755;
    wire tmp4756;
    wire tmp4757;
    wire[7:0] tmp4758;
    wire[7:0] tmp4759;
    wire[8:0] tmp4762;
    wire tmp4763;
    wire tmp4766;
    wire tmp4767;
    wire tmp4768;
    wire tmp4769;
    wire tmp4770;
    wire[6:0] tmp4817;
    wire[6:0] tmp4845;
    wire tmp4874;
    wire[7:0] tmp4876;
    wire tmp4927;
    wire tmp4928;
    wire tmp4992;
    wire tmp5018;
    wire tmp5045;
    wire tmp5069;
    wire tmp5074;
    wire tmp5136;
    wire[8:0] tmp5143;
    wire tmp5144;
    wire tmp5146;
    wire[8:0] tmp5168;
    wire tmp5176;
    wire[6:0] tmp5206;
    wire[7:0] tmp5207;
    wire tmp5226;
    wire tmp5227;
    wire tmp5228;
    wire tmp5229;
    wire tmp5232;
    wire tmp5238;
    wire tmp5259;
    wire[6:0] tmp5287;
    wire tmp5297;
    wire tmp5300;
    wire tmp5306;
    wire tmp5309;
    wire tmp5312;
    wire tmp5313;
    wire tmp5325;
    wire[7:0] tmp5342;
    wire tmp5355;
    wire[8:0] tmp5374;
    wire[8:0] tmp5386;
    wire tmp5387;
    wire tmp5388;
    wire tmp5390;
    wire tmp5418;
    wire tmp5447;
    wire[6:0] tmp5449;
    wire[7:0] tmp5450;
    wire tmp5456;
    wire tmp5462;
    wire[8:0] tmp5467;
    wire tmp5468;
    wire tmp5469;
    wire tmp5470;
    wire tmp5471;
    wire tmp5474;
    wire tmp5475;
    wire tmp5484;
    wire tmp5487;
    wire[8:0] tmp5492;
    wire tmp5493;
    wire tmp5496;
    wire tmp5499;
    wire tmp5500;
    wire tmp5501;
    wire tmp5502;
    wire[7:0] tmp5503;
    wire[7:0] tmp5504;
    wire[8:0] tmp5507;
    wire tmp5508;
    wire tmp5510;
    wire tmp5511;
    wire tmp5512;
    wire tmp5513;
    wire tmp5514;
    wire[8:0] tmp5521;
    wire tmp5525;
    wire tmp5528;
    wire[7:0] tmp5532;
    wire tmp5540;
    wire tmp5541;
    wire[8:0] tmp5546;
    wire tmp5550;
    wire tmp5553;
    wire[7:0] tmp5569;
    wire[7:0] tmp5570;
    wire[8:0] tmp5573;
    wire tmp5574;
    wire tmp5577;
    wire tmp5578;
    wire tmp5579;
    wire tmp5580;
    wire tmp5581;
    wire[6:0] tmp5582;
    wire[7:0] tmp5583;
    wire tmp5595;
    wire[8:0] tmp5600;
    wire tmp5601;
    wire tmp5603;
    wire tmp5604;
    wire tmp5607;
    wire tmp5608;
    wire[8:0] tmp5625;
    wire tmp5626;
    wire tmp5629;
    wire tmp5630;
    wire tmp5632;
    wire tmp5633;
    wire tmp5634;
    wire tmp5635;
    wire[7:0] tmp5636;
    wire[7:0] tmp5637;
    wire[8:0] tmp5640;
    wire tmp5641;
    wire tmp5644;
    wire tmp5645;
    wire tmp5646;
    wire tmp5647;
    wire tmp5648;
    wire tmp5660;
    wire[8:0] tmp5667;
    wire tmp5668;
    wire tmp5674;
    wire[8:0] tmp5680;
    wire[8:0] tmp5692;
    wire tmp5693;
    wire tmp5696;
    wire tmp5699;
    wire tmp5700;
    wire tmp5701;
    wire[8:0] tmp5707;
    wire tmp5708;
    wire tmp5711;
    wire tmp5712;
    wire tmp5713;
    wire tmp5714;
    wire tmp5715;
    wire[6:0] tmp5716;
    wire[7:0] tmp5717;
    wire[8:0] tmp5722;
    wire tmp5723;
    wire tmp5726;
    wire[8:0] tmp5734;
    wire tmp5735;
    wire tmp5737;
    wire tmp5738;
    wire tmp5741;
    wire tmp5742;
    wire tmp5748;
    wire tmp5749;
    wire tmp5751;
    wire[8:0] tmp5759;
    wire tmp5760;
    wire tmp5763;
    wire tmp5764;
    wire tmp5766;
    wire tmp5767;
    wire tmp5768;
    wire tmp5769;
    wire[7:0] tmp5770;
    wire[7:0] tmp5771;
    wire[8:0] tmp5774;
    wire tmp5775;
    wire tmp5778;
    wire tmp5779;
    wire tmp5780;
    wire tmp5781;
    wire tmp5782;
    wire[7:0] tmp5784;
    wire tmp5815;
    wire tmp5831;
    wire tmp5834;
    wire tmp5836;
    wire[8:0] tmp5841;
    wire tmp5842;
    wire tmp5845;
    wire tmp5846;
    wire tmp5847;
    wire tmp5848;
    wire tmp5849;
    wire[6:0] tmp5850;
    wire[7:0] tmp5851;
    wire tmp5863;
    wire[8:0] tmp5868;
    wire tmp5869;
    wire tmp5871;
    wire tmp5872;
    wire tmp5875;
    wire tmp5876;
    wire[8:0] tmp5881;
    wire tmp5882;
    wire tmp5885;
    wire[8:0] tmp5893;
    wire tmp5894;
    wire tmp5897;
    wire tmp5898;
    wire tmp5900;
    wire tmp5901;
    wire tmp5902;
    wire tmp5903;
    wire[7:0] tmp5904;
    wire[7:0] tmp5905;
    wire[8:0] tmp5908;
    wire tmp5909;
    wire tmp5912;
    wire tmp5913;
    wire tmp5914;
    wire tmp5915;
    wire tmp5916;
    wire tmp5942;
    wire[8:0] tmp5960;
    wire tmp5966;
    wire tmp5970;
    wire[7:0] tmp5971;
    wire[8:0] tmp5975;
    wire tmp5976;
    wire tmp5979;
    wire tmp5980;
    wire tmp5981;
    wire tmp5982;
    wire tmp5983;
    wire tmp6058;
    wire[1:0] tmp6067;
    wire[7:0] tmp6074;
    wire[8:0] tmp6079;
    wire tmp6083;
    wire tmp6084;
    wire[8:0] tmp6104;
    wire tmp6105;
    wire tmp6111;
    wire tmp6132;
    wire tmp6138;
    wire tmp6139;
    wire[8:0] tmp6144;
    wire tmp6145;
    wire tmp6148;
    wire tmp6151;
    wire tmp6153;
    wire[7:0] tmp6156;
    wire tmp6205;
    wire[8:0] tmp6210;
    wire[1:0] tmp6211;
    wire[8:0] tmp6213;
    wire[9:0] tmp6221;
    wire[7:0] tmp6222;
    wire tmp6240;
    wire tmp6243;
    wire tmp6244;
    wire tmp6245;
    wire tmp6246;
    wire tmp6247;
    wire tmp6253;
    wire tmp6256;
    wire tmp6259;
    wire tmp6261;
    wire tmp6262;
    wire tmp6274;
    wire[9:0] tmp6279;
    wire tmp6283;
    wire tmp6286;
    wire tmp6287;
    wire[8:0] tmp6292;
    wire tmp6293;
    wire tmp6296;
    wire tmp6297;
    wire tmp6298;
    wire tmp6300;
    wire[7:0] tmp6303;
    wire[7:0] tmp6304;
    wire tmp6355;
    wire[10:0] tmp6368;
    wire[9:0] tmp6369;
    wire[7:0] tmp6370;
    wire[7:0] tmp6384;
    wire tmp6388;
    wire tmp6394;
    wire[8:0] tmp6400;
    wire tmp6401;
    wire tmp6402;
    wire tmp6404;
    wire tmp6407;
    wire tmp6410;
    wire[8:0] tmp6415;
    wire tmp6422;
    wire[9:0] tmp6427;
    wire[8:0] tmp6440;
    wire tmp6444;
    wire tmp6446;
    wire tmp6447;
    wire tmp6449;
    wire tmp6450;
    wire[7:0] tmp6451;
    wire[8:0] tmp6509;
    wire[1:0] tmp6511;
    wire[9:0] tmp6512;
    wire[10:0] tmp6516;
    wire[9:0] tmp6517;
    wire[8:0] tmp6533;
    wire[9:0] tmp6535;
    wire tmp6537;
    wire tmp6538;
    wire tmp6539;
    wire tmp6541;
    wire tmp6542;
    wire tmp6543;
    wire tmp6552;
    wire tmp6555;
    wire tmp6557;
    wire tmp6558;
    wire tmp6570;
    wire[9:0] tmp6575;
    wire tmp6577;
    wire tmp6579;
    wire tmp6583;
    wire[8:0] tmp6588;
    wire tmp6592;
    wire tmp6595;
    wire tmp6597;
    wire tmp6598;
    wire[7:0] tmp6599;
    wire tmp6623;
    wire tmp6651;
    wire tmp6670;
    wire tmp6676;
    wire tmp6725;
    wire[8:0] tmp6734;
    wire[8:0] tmp6735;
    wire[8:0] tmp6744;
    wire[8:0] tmp6746;
    wire[8:0] tmp6747;
    wire[9:0] tmp6750;
    wire tmp6751;
    wire tmp6752;
    wire tmp6753;
    wire tmp6754;
    wire tmp6755;
    wire tmp6756;
    wire tmp6757;
    wire tmp6759;
    wire[8:0] tmp6763;
    wire[8:0] tmp6766;
    wire[8:0] tmp6769;
    wire tmp6771;
    wire[8:0] tmp6780;
    wire[8:0] tmp6781;
    wire[9:0] tmp6784;
    wire tmp6785;
    wire tmp6786;
    wire tmp6787;
    wire tmp6788;
    wire tmp6789;
    wire tmp6790;
    wire tmp6791;
    wire tmp6792;
    wire[8:0] tmp6803;
    wire tmp6807;
    wire[8:0] tmp6813;
    wire[9:0] tmp6819;
    wire tmp6820;
    wire tmp6821;
    wire tmp6822;
    wire tmp6823;
    wire tmp6825;
    wire tmp6826;
    wire tmp6827;
    wire tmp6829;
    wire tmp6830;
    wire[8:0] tmp6838;
    wire[8:0] tmp6839;
    wire tmp6841;
    wire[8:0] tmp6845;
    wire[8:0] tmp6848;
    wire[9:0] tmp6854;
    wire tmp6855;
    wire tmp6856;
    wire tmp6857;
    wire tmp6858;
    wire tmp6859;
    wire tmp6861;
    wire tmp6862;
    wire tmp6958;
    wire tmp6972;
    wire[7:0] tmp7035;
    wire tmp7036;
    wire[8:0] tmp7038;
    wire tmp7040;
    wire tmp7041;
    wire[9:0] tmp7053;
    wire tmp7054;
    wire tmp7055;
    wire tmp7056;
    wire tmp7057;
    wire tmp7060;
    wire tmp7061;
    wire tmp7062;
    wire tmp7063;
    wire[8:0] tmp7074;
    wire[7:0] tmp7076;
    wire tmp7077;
    wire[8:0] tmp7079;
    wire[8:0] tmp7088;
    wire[9:0] tmp7094;
    wire tmp7095;
    wire tmp7096;
    wire tmp7097;
    wire tmp7098;
    wire tmp7101;
    wire tmp7102;
    wire tmp7103;
    wire tmp7104;
    wire tmp7106;
    wire[8:0] tmp7116;
    wire[7:0] tmp7117;
    wire tmp7118;
    wire[8:0] tmp7120;
    wire tmp7121;
    wire tmp7122;
    wire[8:0] tmp7131;
    wire[8:0] tmp7132;
    wire[9:0] tmp7135;
    wire tmp7136;
    wire tmp7137;
    wire tmp7138;
    wire tmp7139;
    wire tmp7140;
    wire tmp7142;
    wire tmp7143;
    wire tmp7144;
    wire tmp7145;
    wire[7:0] tmp7158;
    wire tmp7159;
    wire[8:0] tmp7161;
    wire tmp7162;
    wire[8:0] tmp7172;
    wire[8:0] tmp7173;
    wire[9:0] tmp7176;
    wire tmp7177;
    wire tmp7178;
    wire tmp7179;
    wire tmp7180;
    wire tmp7182;
    wire tmp7183;
    wire tmp7184;
    wire tmp7185;
    wire tmp7186;
    wire[6:0] tmp7223;
    wire tmp7224;
    wire[7:0] tmp7226;
    wire tmp7242;
    wire tmp7243;
    wire tmp7244;
    wire[6:0] tmp7246;
    wire tmp7247;
    wire[7:0] tmp7249;
    wire tmp7268;
    wire[6:0] tmp7269;
    wire tmp7270;
    wire[7:0] tmp7272;
    wire[6:0] tmp7292;
    wire tmp7293;
    wire[7:0] tmp7295;
    wire[7:0] tmp7316;
    wire[8:0] tmp7321;
    wire tmp7325;
    wire tmp7327;
    wire tmp7341;
    wire[8:0] tmp7358;
    wire tmp7362;
    wire tmp7366;
    wire tmp7368;
    wire[7:0] tmp7370;
    wire tmp7383;
    wire[6:0] tmp7391;
    wire[7:0] tmp7392;
    wire tmp7404;
    wire[8:0] tmp7409;
    wire tmp7411;
    wire tmp7412;
    wire tmp7413;
    wire tmp7416;
    wire tmp7417;
    wire[8:0] tmp7422;
    wire[8:0] tmp7434;
    wire tmp7435;
    wire tmp7438;
    wire tmp7441;
    wire tmp7442;
    wire tmp7443;
    wire[7:0] tmp7445;
    wire[7:0] tmp7446;
    wire tmp7466;
    wire[6:0] tmp7467;
    wire[7:0] tmp7468;
    wire tmp7474;
    wire tmp7486;
    wire tmp7487;
    wire tmp7488;
    wire tmp7493;
    wire tmp7502;
    wire tmp7517;
    wire tmp7518;
    wire[6:0] tmp7543;
    wire[7:0] tmp7544;
    wire tmp7556;
    wire[8:0] tmp7561;
    wire tmp7562;
    wire tmp7563;
    wire tmp7565;
    wire tmp7568;
    wire tmp7569;
    wire[8:0] tmp7586;
    wire tmp7587;
    wire tmp7590;
    wire tmp7592;
    wire tmp7593;
    wire tmp7594;
    wire tmp7595;
    wire tmp7596;
    wire[7:0] tmp7597;
    wire[7:0] tmp7598;
    wire tmp7636;
    wire tmp7637;
    wire tmp7644;
    wire[7:0] tmp7689;
    wire[7:0] tmp7690;
    wire[7:0] tmp7691;
    wire[7:0] tmp7692;
    wire[7:0] tmp7693;
    wire[7:0] tmp7694;
    wire[7:0] tmp7695;
    wire[7:0] tmp7696;
    wire[7:0] tmp7697;
    wire[7:0] tmp7698;
    wire[7:0] tmp7699;
    wire[7:0] tmp7700;
    wire[7:0] tmp7701;
    wire[7:0] tmp7702;
    wire[7:0] tmp7703;
    wire[7:0] tmp7704;
    wire[7:0] tmp7705;
    wire[7:0] tmp7706;
    wire[7:0] tmp7707;
    wire[7:0] tmp7708;
    wire[7:0] tmp7709;
    wire[7:0] tmp7710;
    wire[7:0] tmp7711;
    wire[7:0] tmp7712;
    wire[7:0] tmp7713;
    wire[7:0] tmp7714;
    wire[7:0] tmp7715;
    wire[7:0] tmp7716;
    wire[7:0] tmp7717;
    wire[7:0] tmp7718;
    wire[7:0] tmp7719;
    wire[7:0] tmp7720;
    wire[7:0] tmp7721;
    wire[7:0] tmp7722;
    wire[7:0] tmp7723;
    wire[7:0] tmp7724;
    wire[7:0] tmp7725;
    wire[7:0] tmp7726;
    wire[7:0] tmp7727;
    wire[7:0] tmp7728;
    wire[7:0] tmp7729;
    wire[7:0] tmp7730;
    wire[7:0] tmp7731;
    wire[7:0] tmp7732;
    wire[7:0] tmp7733;
    wire[7:0] tmp7734;
    wire[7:0] tmp7735;
    wire[7:0] tmp7736;
    wire[7:0] tmp7737;
    wire[7:0] tmp7738;
    wire[7:0] tmp7739;
    wire[7:0] tmp7740;
    wire[7:0] tmp7741;
    wire[7:0] tmp7742;
    wire[7:0] tmp7743;
    wire[7:0] tmp7744;
    wire[7:0] tmp7745;
    wire[7:0] tmp7746;
    wire[7:0] tmp7747;
    wire[7:0] tmp7748;
    wire[7:0] tmp7749;
    wire[7:0] tmp7750;
    wire[7:0] tmp7751;
    wire[7:0] tmp7752;
    wire[7:0] tmp7753;
    wire[7:0] tmp7754;
    wire[7:0] tmp7755;
    wire[7:0] tmp7756;
    wire[7:0] tmp7757;
    wire[7:0] tmp7758;
    wire[7:0] tmp7759;
    wire[7:0] tmp7760;
    wire[7:0] tmp7761;
    wire[7:0] tmp7762;
    wire[7:0] tmp7763;
    wire[7:0] tmp7764;
    wire[7:0] tmp7765;
    wire[7:0] tmp7766;
    wire[7:0] tmp7767;
    wire[7:0] tmp7768;
    wire[7:0] tmp7769;
    wire[7:0] tmp7770;
    wire[7:0] tmp7771;
    wire[7:0] tmp7772;
    wire[7:0] tmp7773;
    wire[7:0] tmp7774;
    wire[7:0] tmp7775;
    wire[7:0] tmp7776;
    wire[7:0] tmp7777;
    wire[7:0] tmp7778;
    wire[7:0] tmp7779;
    wire[7:0] tmp7780;
    wire[7:0] tmp7781;
    wire[7:0] tmp7782;
    wire[7:0] tmp7783;
    wire[7:0] tmp7784;
    wire[7:0] tmp7785;
    wire[7:0] tmp7786;
    wire[7:0] tmp7787;
    wire[7:0] tmp7788;
    wire[7:0] tmp7789;
    wire[7:0] tmp7790;
    wire[7:0] tmp7791;
    wire[7:0] tmp7792;
    wire[7:0] tmp7793;
    wire[7:0] tmp7794;
    wire[7:0] tmp7795;
    wire[7:0] tmp7796;
    wire[7:0] tmp7797;
    wire[7:0] tmp7798;
    wire[7:0] tmp7799;
    wire[7:0] tmp7800;
    wire[7:0] tmp7801;
    wire[7:0] tmp7802;
    wire[7:0] tmp7803;
    wire[7:0] tmp7804;
    wire[7:0] tmp7805;
    wire[7:0] tmp7806;
    wire[7:0] tmp7807;
    wire[7:0] tmp7808;
    wire[7:0] tmp7809;
    wire[7:0] tmp7810;
    wire[7:0] tmp7811;
    wire[7:0] tmp7812;
    wire[7:0] tmp7813;
    wire[7:0] tmp7814;
    wire[7:0] tmp7815;
    wire[7:0] tmp7816;
    wire[7:0] tmp7817;
    wire[7:0] tmp7818;
    wire[7:0] tmp7819;
    wire[7:0] tmp7820;
    wire[7:0] tmp7821;
    wire[7:0] tmp7822;
    wire[7:0] tmp7823;
    wire[7:0] tmp7824;
    wire[7:0] tmp7825;
    wire[7:0] tmp7826;
    wire[7:0] tmp7827;
    wire[7:0] tmp7828;
    wire tmp7829;
    wire tmp7830;
    wire tmp7831;
    wire tmp7832;
    wire tmp7833;
    wire tmp7834;
    wire tmp7835;
    wire tmp7836;
    wire tmp7837;
    wire tmp7838;
    wire tmp7839;
    wire tmp7840;
    wire tmp7841;
    wire tmp7842;
    wire tmp7843;
    wire tmp7844;
    wire tmp7845;
    wire tmp7846;
    wire tmp7847;
    wire tmp7848;
    wire tmp7849;
    wire[7:0] tmp7852;
    wire[7:0] tmp7853;
    wire[7:0] tmp7856;
    wire[7:0] tmp7857;
    wire[7:0] tmp7860;
    wire[7:0] tmp7861;
    wire[7:0] tmp7864;
    wire[7:0] tmp7865;
    wire[7:0] tmp7868;
    wire[7:0] tmp7869;
    wire[7:0] tmp7872;
    wire[7:0] tmp7873;
    wire[7:0] tmp7876;
    wire[7:0] tmp7877;
    wire[7:0] tmp7880;
    wire[7:0] tmp7881;
    wire[3:0] tmp7882;
    wire[3:0] tmp7883;
    wire[3:0] tmp7884;
    wire[3:0] tmp7885;
    wire[3:0] tmp7886;
    wire[3:0] tmp7887;
    wire[3:0] tmp7888;
    wire[3:0] tmp7889;
    wire[3:0] tmp7890;
    wire[3:0] tmp7891;
    wire[3:0] tmp7892;
    wire[3:0] tmp7893;
    wire[3:0] tmp7894;
    wire tmp7902;
    wire[3:0] tmp7904;
    wire tmp7905;
    wire tmp7906;
    wire[3:0] tmp7908;
    wire tmp7909;
    wire tmp7910;
    wire tmp7912;
    wire tmp7915;
    wire[3:0] tmp7917;
    wire tmp7918;
    wire tmp7919;
    wire tmp7923;
    wire tmp7926;
    wire tmp7927;
    wire tmp7929;
    wire tmp7930;
    wire tmp7933;
    wire tmp7934;
    wire tmp7938;
    wire tmp7939;
    wire tmp7940;
    wire[2:0] tmp7941;
    wire[3:0] tmp7942;
    wire[3:0] tmp7943;
    wire[3:0] tmp7944;
    wire[4:0] tmp7945;
    wire[5:0] tmp7946;
    wire[4:0] tmp7947;
    wire tmp7949;
    wire tmp7950;
    wire tmp7953;
    wire tmp7954;
    wire tmp7956;
    wire tmp7959;
    wire tmp7961;
    wire tmp7962;
    wire tmp7963;
    wire tmp7964;
    wire tmp7967;
    wire tmp7972;
    wire tmp7973;
    wire tmp7974;
    wire[4:0] tmp7975;
    wire[3:0] tmp7976;
    wire[3:0] tmp7977;
    wire[3:0] tmp7978;
    wire[3:0] tmp7979;

    initial begin
        mem_0[0]=3'h4;
        mem_0[1]=3'h1;
        mem_0[2]=3'h2;
        mem_0[3]=3'h3;
        mem_0[4]=3'h1;
        mem_0[5]=3'h2;
        mem_0[6]=3'h3;
        mem_0[7]=3'h1;
        mem_0[8]=3'h2;
        mem_0[9]=3'h3;
        mem_0[10]=3'h1;
        mem_0[11]=3'h2;
        mem_0[12]=3'h3;
        mem_0[13]=3'h1;
        mem_0[14]=3'h2;
        mem_0[15]=3'h3;
        mem_0[16]=3'h1;
        mem_0[17]=3'h2;
        mem_0[18]=3'h3;
        mem_0[19]=3'h1;
        mem_0[20]=3'h2;
        mem_0[21]=3'h3;
        mem_0[22]=3'h1;
        mem_0[23]=3'h2;
        mem_0[24]=3'h3;
        mem_0[25]=3'h1;
        mem_0[26]=3'h2;
        mem_0[27]=3'h3;
        mem_0[28]=3'h1;
        mem_0[29]=3'h2;
        mem_0[30]=3'h3;
        mem_0[31]=3'h1;
    end

    initial begin
        mem_1[0]=4'h0;
        mem_1[1]=4'h4;
        mem_1[2]=4'h4;
        mem_1[3]=4'h4;
        mem_1[4]=4'hf;
        mem_1[5]=4'hf;
        mem_1[6]=4'hf;
        mem_1[7]=4'h0;
        mem_1[8]=4'h0;
        mem_1[9]=4'h0;
        mem_1[10]=4'h0;
        mem_1[11]=4'h0;
        mem_1[12]=4'h0;
        mem_1[13]=4'h0;
        mem_1[14]=4'h0;
        mem_1[15]=4'h0;
        mem_1[16]=4'h0;
        mem_1[17]=4'h0;
        mem_1[18]=4'h0;
        mem_1[19]=4'h0;
        mem_1[20]=4'h0;
        mem_1[21]=4'h0;
        mem_1[22]=4'h0;
        mem_1[23]=4'h0;
        mem_1[24]=4'h0;
        mem_1[25]=4'h0;
        mem_1[26]=4'h0;
        mem_1[27]=4'h0;
        mem_1[28]=4'h0;
        mem_1[29]=4'h0;
        mem_1[30]=4'h0;
        mem_1[31]=4'h0;
    end

    initial begin
        mem_2[0]=4'h0;
        mem_2[1]=4'h1;
        mem_2[2]=4'h1;
        mem_2[3]=4'h1;
        mem_2[4]=4'h4;
        mem_2[5]=4'h4;
        mem_2[6]=4'h4;
        mem_2[7]=4'hf;
        mem_2[8]=4'hf;
        mem_2[9]=4'hf;
        mem_2[10]=4'h0;
        mem_2[11]=4'h0;
        mem_2[12]=4'h0;
        mem_2[13]=4'h0;
        mem_2[14]=4'h0;
        mem_2[15]=4'h0;
        mem_2[16]=4'h0;
        mem_2[17]=4'h0;
        mem_2[18]=4'h0;
        mem_2[19]=4'h0;
        mem_2[20]=4'h0;
        mem_2[21]=4'h0;
        mem_2[22]=4'h0;
        mem_2[23]=4'h0;
        mem_2[24]=4'h0;
        mem_2[25]=4'h0;
        mem_2[26]=4'h0;
        mem_2[27]=4'h0;
        mem_2[28]=4'h0;
        mem_2[29]=4'h0;
        mem_2[30]=4'h0;
        mem_2[31]=4'h0;
    end

    // Combinational
    assign _ver_out_tmp_0 = 128;
    assign _ver_out_tmp_1 = 128;
    assign _ver_out_tmp_2 = 128;
    assign _ver_out_tmp_3 = 128;
    assign _ver_out_tmp_4 = 128;
    assign _ver_out_tmp_5 = 128;
    assign _ver_out_tmp_6 = 128;
    assign _ver_out_tmp_7 = 128;
    assign _ver_out_tmp_8 = 128;
    assign _ver_out_tmp_9 = 128;
    assign _ver_out_tmp_10 = 128;
    assign _ver_out_tmp_11 = 128;
    assign _ver_out_tmp_12 = 128;
    assign _ver_out_tmp_13 = 128;
    assign _ver_out_tmp_14 = 128;
    assign _ver_out_tmp_15 = 128;
    assign _ver_out_tmp_16 = 128;
    assign _ver_out_tmp_17 = 128;
    assign _ver_out_tmp_18 = 128;
    assign _ver_out_tmp_19 = 128;
    assign _ver_out_tmp_20 = 128;
    assign _ver_out_tmp_21 = 128;
    assign _ver_out_tmp_22 = 128;
    assign _ver_out_tmp_23 = 128;
    assign _ver_out_tmp_24 = 128;
    assign _ver_out_tmp_25 = 128;
    assign _ver_out_tmp_26 = 128;
    assign _ver_out_tmp_27 = 128;
    assign _ver_out_tmp_28 = 128;
    assign _ver_out_tmp_29 = 128;
    assign _ver_out_tmp_30 = 128;
    assign _ver_out_tmp_31 = 128;
    assign _ver_out_tmp_32 = 128;
    assign _ver_out_tmp_33 = 128;
    assign _ver_out_tmp_34 = 128;
    assign _ver_out_tmp_35 = 128;
    assign _ver_out_tmp_36 = 128;
    assign _ver_out_tmp_37 = 128;
    assign _ver_out_tmp_38 = 128;
    assign _ver_out_tmp_39 = 128;
    assign _ver_out_tmp_40 = 128;
    assign _ver_out_tmp_41 = 128;
    assign _ver_out_tmp_42 = 128;
    assign _ver_out_tmp_43 = 128;
    assign _ver_out_tmp_44 = 128;
    assign _ver_out_tmp_45 = 128;
    assign _ver_out_tmp_46 = 128;
    assign _ver_out_tmp_47 = 128;
    assign _ver_out_tmp_48 = 128;
    assign _ver_out_tmp_49 = 128;
    assign _ver_out_tmp_50 = 128;
    assign _ver_out_tmp_51 = 128;
    assign _ver_out_tmp_52 = 128;
    assign _ver_out_tmp_53 = 128;
    assign _ver_out_tmp_54 = 128;
    assign _ver_out_tmp_55 = 128;
    assign _ver_out_tmp_56 = 128;
    assign _ver_out_tmp_57 = 128;
    assign _ver_out_tmp_58 = 128;
    assign _ver_out_tmp_59 = 128;
    assign _ver_out_tmp_60 = 128;
    assign _ver_out_tmp_61 = 128;
    assign _ver_out_tmp_62 = 128;
    assign _ver_out_tmp_63 = 128;
    assign _ver_out_tmp_64 = 128;
    assign _ver_out_tmp_65 = 128;
    assign _ver_out_tmp_66 = 128;
    assign _ver_out_tmp_67 = 128;
    assign _ver_out_tmp_68 = 128;
    assign _ver_out_tmp_69 = 128;
    assign _ver_out_tmp_70 = 128;
    assign _ver_out_tmp_71 = 128;
    assign _ver_out_tmp_72 = 128;
    assign _ver_out_tmp_73 = 128;
    assign _ver_out_tmp_74 = 128;
    assign _ver_out_tmp_75 = 128;
    assign _ver_out_tmp_76 = 128;
    assign _ver_out_tmp_77 = 128;
    assign _ver_out_tmp_78 = 128;
    assign _ver_out_tmp_79 = 128;
    assign _ver_out_tmp_80 = 128;
    assign _ver_out_tmp_81 = 128;
    assign _ver_out_tmp_82 = 128;
    assign _ver_out_tmp_83 = 128;
    assign _ver_out_tmp_84 = 128;
    assign _ver_out_tmp_85 = 128;
    assign _ver_out_tmp_86 = 128;
    assign _ver_out_tmp_87 = 128;
    assign _ver_out_tmp_88 = 128;
    assign _ver_out_tmp_89 = 128;
    assign _ver_out_tmp_90 = 128;
    assign _ver_out_tmp_91 = 128;
    assign const_1_1 = 1;
    assign const_2_0 = 0;
    assign const_3_0 = 0;
    assign const_4_0 = 0;
    assign const_5_4 = 4;
    assign const_6_0 = 0;
    assign const_7_2 = 2;
    assign const_8_1 = 1;
    assign const_9_0 = 0;
    assign const_10_0 = 0;
    assign const_11_0 = 0;
    assign const_12_0 = 0;
    assign const_13_1 = 1;
    assign const_14_0 = 0;
    assign const_15_1 = 1;
    assign const_16_0 = 0;
    assign const_17_0 = 0;
    assign const_18_0 = 0;
    assign const_19_15 = 15;
    assign const_20_1 = 1;
    assign const_21_0 = 0;
    assign const_22_2 = 2;
    assign const_23_0 = 0;
    assign const_24_3 = 3;
    assign const_25_0 = 0;
    assign const_26_0 = 0;
    assign const_27_0 = 0;
    assign const_28_0 = 0;
    assign const_29_0 = 0;
    assign const_30_0 = 0;
    assign const_31_127 = 127;
    assign const_33_0 = 0;
    assign const_34_0 = 0;
    assign const_35_0 = 0;
    assign const_36_0 = 0;
    assign const_37_0 = 0;
    assign const_38_127 = 127;
    assign const_40_0 = 0;
    assign const_41_0 = 0;
    assign const_42_0 = 0;
    assign const_43_0 = 0;
    assign const_44_0 = 0;
    assign const_45_127 = 127;
    assign const_47_0 = 0;
    assign const_48_0 = 0;
    assign const_49_0 = 0;
    assign const_50_0 = 0;
    assign const_51_0 = 0;
    assign const_52_127 = 127;
    assign const_54_6 = 6;
    assign const_55_0 = 0;
    assign const_56_7 = 7;
    assign const_57_0 = 0;
    assign const_58_4 = 4;
    assign const_59_0 = 0;
    assign const_60_5 = 5;
    assign const_61_0 = 0;
    assign const_62_0 = 0;
    assign const_63_0 = 0;
    assign const_64_0 = 0;
    assign const_65_0 = 0;
    assign const_66_0 = 0;
    assign const_67_0 = 0;
    assign const_68_127 = 127;
    assign const_70_0 = 0;
    assign const_71_0 = 0;
    assign const_72_0 = 0;
    assign const_73_0 = 0;
    assign const_74_0 = 0;
    assign const_75_0 = 0;
    assign const_76_127 = 127;
    assign const_78_0 = 0;
    assign const_79_0 = 0;
    assign const_80_0 = 0;
    assign const_81_0 = 0;
    assign const_82_0 = 0;
    assign const_83_0 = 0;
    assign const_84_127 = 127;
    assign const_86_0 = 0;
    assign const_87_0 = 0;
    assign const_88_0 = 0;
    assign const_89_0 = 0;
    assign const_90_0 = 0;
    assign const_91_0 = 0;
    assign const_92_127 = 127;
    assign const_94_8 = 8;
    assign const_96_0 = 0;
    assign const_97_0 = 0;
    assign const_98_127 = 127;
    assign const_99_0 = 0;
    assign const_101_0 = 0;
    assign const_102_0 = 0;
    assign const_103_127 = 127;
    assign const_104_0 = 0;
    assign const_106_0 = 0;
    assign const_107_0 = 0;
    assign const_108_127 = 127;
    assign const_109_0 = 0;
    assign const_111_0 = 0;
    assign const_112_0 = 0;
    assign const_113_127 = 127;
    assign const_114_0 = 0;
    assign const_115_2 = 2;
    assign const_116_0 = 0;
    assign const_117_0 = 0;
    assign const_118_0 = 0;
    assign const_119_15 = 15;
    assign const_120_1 = 1;
    assign const_121_0 = 0;
    assign const_122_2 = 2;
    assign const_123_0 = 0;
    assign const_124_3 = 3;
    assign const_125_0 = 0;
    assign const_126_0 = 0;
    assign const_127_0 = 0;
    assign const_128_0 = 0;
    assign const_129_0 = 0;
    assign const_130_0 = 0;
    assign const_131_127 = 127;
    assign const_133_0 = 0;
    assign const_134_0 = 0;
    assign const_135_0 = 0;
    assign const_136_0 = 0;
    assign const_137_0 = 0;
    assign const_138_127 = 127;
    assign const_140_0 = 0;
    assign const_141_0 = 0;
    assign const_142_0 = 0;
    assign const_143_0 = 0;
    assign const_144_0 = 0;
    assign const_145_127 = 127;
    assign const_147_0 = 0;
    assign const_148_0 = 0;
    assign const_149_0 = 0;
    assign const_150_0 = 0;
    assign const_151_0 = 0;
    assign const_152_127 = 127;
    assign const_154_6 = 6;
    assign const_155_0 = 0;
    assign const_156_7 = 7;
    assign const_157_0 = 0;
    assign const_158_4 = 4;
    assign const_159_0 = 0;
    assign const_160_5 = 5;
    assign const_161_0 = 0;
    assign const_162_0 = 0;
    assign const_163_0 = 0;
    assign const_164_0 = 0;
    assign const_165_0 = 0;
    assign const_166_0 = 0;
    assign const_167_0 = 0;
    assign const_168_127 = 127;
    assign const_170_0 = 0;
    assign const_171_0 = 0;
    assign const_172_0 = 0;
    assign const_173_0 = 0;
    assign const_174_0 = 0;
    assign const_175_0 = 0;
    assign const_176_127 = 127;
    assign const_178_0 = 0;
    assign const_179_0 = 0;
    assign const_180_0 = 0;
    assign const_181_0 = 0;
    assign const_182_0 = 0;
    assign const_183_0 = 0;
    assign const_184_127 = 127;
    assign const_186_0 = 0;
    assign const_187_0 = 0;
    assign const_188_0 = 0;
    assign const_189_0 = 0;
    assign const_190_0 = 0;
    assign const_191_0 = 0;
    assign const_192_127 = 127;
    assign const_194_8 = 8;
    assign const_196_0 = 0;
    assign const_197_0 = 0;
    assign const_198_127 = 127;
    assign const_199_0 = 0;
    assign const_201_0 = 0;
    assign const_202_0 = 0;
    assign const_203_127 = 127;
    assign const_204_0 = 0;
    assign const_206_0 = 0;
    assign const_207_0 = 0;
    assign const_208_127 = 127;
    assign const_209_0 = 0;
    assign const_211_0 = 0;
    assign const_212_0 = 0;
    assign const_213_127 = 127;
    assign const_214_0 = 0;
    assign const_215_3 = 3;
    assign const_216_0 = 0;
    assign const_217_0 = 0;
    assign const_218_0 = 0;
    assign const_219_0 = 0;
    assign const_220_0 = 0;
    assign const_221_0 = 0;
    assign const_222_0 = 0;
    assign const_223_0 = 0;
    assign const_224_0 = 0;
    assign const_225_0 = 0;
    assign const_226_0 = 0;
    assign const_227_0 = 0;
    assign const_228_0 = 0;
    assign const_229_0 = 0;
    assign const_230_0 = 0;
    assign const_231_0 = 0;
    assign const_232_0 = 0;
    assign const_233_0 = 0;
    assign const_234_0 = 0;
    assign const_235_0 = 0;
    assign const_236_0 = 0;
    assign const_237_0 = 0;
    assign const_238_0 = 0;
    assign const_240_0 = 0;
    assign const_241_0 = 0;
    assign const_242_127 = 127;
    assign const_243_0 = 0;
    assign const_245_0 = 0;
    assign const_246_0 = 0;
    assign const_247_127 = 127;
    assign const_248_0 = 0;
    assign const_250_0 = 0;
    assign const_251_0 = 0;
    assign const_252_127 = 127;
    assign const_253_0 = 0;
    assign const_255_0 = 0;
    assign const_256_0 = 0;
    assign const_257_127 = 127;
    assign const_258_0 = 0;
    assign const_260_0 = 0;
    assign const_261_0 = 0;
    assign const_262_127 = 127;
    assign const_263_0 = 0;
    assign const_265_0 = 0;
    assign const_266_0 = 0;
    assign const_267_127 = 127;
    assign const_268_0 = 0;
    assign const_270_0 = 0;
    assign const_271_0 = 0;
    assign const_272_127 = 127;
    assign const_273_0 = 0;
    assign const_275_0 = 0;
    assign const_276_0 = 0;
    assign const_277_127 = 127;
    assign const_278_0 = 0;
    assign const_279_0 = 0;
    assign const_280_0 = 0;
    assign const_281_0 = 0;
    assign const_282_0 = 0;
    assign const_283_0 = 0;
    assign const_284_0 = 0;
    assign const_285_0 = 0;
    assign const_286_0 = 0;
    assign const_287_0 = 0;
    assign const_288_0 = 0;
    assign const_289_15 = 15;
    assign const_290_0 = 0;
    assign const_291_0 = 0;
    assign const_292_0 = 0;
    assign const_293_8 = 8;
    assign const_294_0 = 0;
    assign const_296_0 = 0;
    assign const_297_0 = 0;
    assign const_298_127 = 127;
    assign const_299_0 = 0;
    assign const_301_0 = 0;
    assign const_302_0 = 0;
    assign const_303_127 = 127;
    assign const_304_0 = 0;
    assign const_306_0 = 0;
    assign const_307_0 = 0;
    assign const_308_127 = 127;
    assign const_309_0 = 0;
    assign const_311_0 = 0;
    assign const_312_0 = 0;
    assign const_313_127 = 127;
    assign const_314_0 = 0;
    assign const_315_1 = 1;
    assign const_316_0 = 0;
    assign const_317_0 = 0;
    assign const_318_0 = 0;
    assign const_319_0 = 0;
    assign const_320_0 = 0;
    assign const_321_0 = 0;
    assign const_322_127 = 127;
    assign const_324_0 = 0;
    assign const_325_0 = 0;
    assign const_326_0 = 0;
    assign const_327_0 = 0;
    assign const_328_0 = 0;
    assign const_329_127 = 127;
    assign const_331_0 = 0;
    assign const_332_0 = 0;
    assign const_333_0 = 0;
    assign const_334_0 = 0;
    assign const_335_0 = 0;
    assign const_336_127 = 127;
    assign const_338_0 = 0;
    assign const_339_0 = 0;
    assign const_340_0 = 0;
    assign const_341_0 = 0;
    assign const_342_0 = 0;
    assign const_343_127 = 127;
    assign const_345_4 = 4;
    assign const_346_0 = 0;
    assign const_348_0 = 0;
    assign const_349_0 = 0;
    assign const_350_127 = 127;
    assign const_351_0 = 0;
    assign const_352_0 = 0;
    assign const_353_0 = 0;
    assign const_354_0 = 0;
    assign const_355_0 = 0;
    assign const_356_0 = 0;
    assign const_357_0 = 0;
    assign const_358_127 = 127;
    assign const_361_0 = 0;
    assign const_362_0 = 0;
    assign const_363_127 = 127;
    assign const_364_0 = 0;
    assign const_365_0 = 0;
    assign const_366_0 = 0;
    assign const_367_0 = 0;
    assign const_368_0 = 0;
    assign const_369_0 = 0;
    assign const_370_0 = 0;
    assign const_371_127 = 127;
    assign const_374_0 = 0;
    assign const_375_0 = 0;
    assign const_376_127 = 127;
    assign const_377_0 = 0;
    assign const_378_0 = 0;
    assign const_379_0 = 0;
    assign const_380_0 = 0;
    assign const_381_0 = 0;
    assign const_382_0 = 0;
    assign const_383_0 = 0;
    assign const_384_127 = 127;
    assign const_387_0 = 0;
    assign const_388_0 = 0;
    assign const_389_127 = 127;
    assign const_390_0 = 0;
    assign const_391_0 = 0;
    assign const_392_0 = 0;
    assign const_393_0 = 0;
    assign const_394_0 = 0;
    assign const_395_0 = 0;
    assign const_396_0 = 0;
    assign const_397_127 = 127;
    assign const_399_6 = 6;
    assign const_400_0 = 0;
    assign const_401_0 = 0;
    assign const_402_0 = 0;
    assign const_403_0 = 0;
    assign const_404_0 = 0;
    assign const_405_0 = 0;
    assign const_406_127 = 127;
    assign const_408_0 = 0;
    assign const_409_0 = 0;
    assign const_410_0 = 0;
    assign const_411_0 = 0;
    assign const_412_0 = 0;
    assign const_413_127 = 127;
    assign const_415_0 = 0;
    assign const_416_0 = 0;
    assign const_417_0 = 0;
    assign const_418_0 = 0;
    assign const_419_0 = 0;
    assign const_420_127 = 127;
    assign const_422_0 = 0;
    assign const_423_0 = 0;
    assign const_424_0 = 0;
    assign const_425_0 = 0;
    assign const_426_0 = 0;
    assign const_427_127 = 127;
    assign const_429_2 = 2;
    assign const_430_0 = 0;
    assign const_431_0 = 0;
    assign const_432_0 = 0;
    assign const_433_0 = 0;
    assign const_434_0 = 0;
    assign const_435_0 = 0;
    assign const_436_127 = 127;
    assign const_438_0 = 0;
    assign const_439_0 = 0;
    assign const_440_0 = 0;
    assign const_441_0 = 0;
    assign const_442_0 = 0;
    assign const_443_127 = 127;
    assign const_445_0 = 0;
    assign const_446_0 = 0;
    assign const_447_0 = 0;
    assign const_448_0 = 0;
    assign const_449_0 = 0;
    assign const_450_127 = 127;
    assign const_452_0 = 0;
    assign const_453_0 = 0;
    assign const_454_0 = 0;
    assign const_455_0 = 0;
    assign const_456_0 = 0;
    assign const_457_127 = 127;
    assign const_459_0 = 0;
    assign const_460_0 = 0;
    assign const_461_0 = 0;
    assign const_462_0 = 0;
    assign const_463_0 = 0;
    assign const_464_127 = 127;
    assign const_466_0 = 0;
    assign const_467_0 = 0;
    assign const_468_0 = 0;
    assign const_469_0 = 0;
    assign const_470_0 = 0;
    assign const_471_127 = 127;
    assign const_473_0 = 0;
    assign const_474_0 = 0;
    assign const_475_0 = 0;
    assign const_476_0 = 0;
    assign const_477_0 = 0;
    assign const_478_127 = 127;
    assign const_480_0 = 0;
    assign const_481_0 = 0;
    assign const_482_0 = 0;
    assign const_483_0 = 0;
    assign const_484_0 = 0;
    assign const_485_127 = 127;
    assign const_487_0 = 0;
    assign const_488_0 = 0;
    assign const_489_0 = 0;
    assign const_490_0 = 0;
    assign const_491_0 = 0;
    assign const_492_127 = 127;
    assign const_494_0 = 0;
    assign const_495_0 = 0;
    assign const_496_0 = 0;
    assign const_497_0 = 0;
    assign const_498_0 = 0;
    assign const_499_127 = 127;
    assign const_501_0 = 0;
    assign const_502_0 = 0;
    assign const_503_0 = 0;
    assign const_504_0 = 0;
    assign const_505_0 = 0;
    assign const_506_127 = 127;
    assign const_508_0 = 0;
    assign const_509_0 = 0;
    assign const_510_0 = 0;
    assign const_511_0 = 0;
    assign const_512_0 = 0;
    assign const_513_127 = 127;
    assign const_515_5 = 5;
    assign const_516_1 = 1;
    assign const_518_0 = 0;
    assign const_519_0 = 0;
    assign const_520_127 = 127;
    assign const_521_0 = 0;
    assign const_522_0 = 0;
    assign const_523_0 = 0;
    assign const_524_0 = 0;
    assign const_525_0 = 0;
    assign const_526_0 = 0;
    assign const_527_0 = 0;
    assign const_528_127 = 127;
    assign const_531_0 = 0;
    assign const_532_0 = 0;
    assign const_533_127 = 127;
    assign const_534_0 = 0;
    assign const_535_0 = 0;
    assign const_536_0 = 0;
    assign const_537_0 = 0;
    assign const_538_0 = 0;
    assign const_539_0 = 0;
    assign const_540_0 = 0;
    assign const_541_127 = 127;
    assign const_544_0 = 0;
    assign const_545_0 = 0;
    assign const_546_127 = 127;
    assign const_547_0 = 0;
    assign const_548_0 = 0;
    assign const_549_0 = 0;
    assign const_550_0 = 0;
    assign const_551_0 = 0;
    assign const_552_0 = 0;
    assign const_553_0 = 0;
    assign const_554_127 = 127;
    assign const_557_0 = 0;
    assign const_558_0 = 0;
    assign const_559_127 = 127;
    assign const_560_0 = 0;
    assign const_561_0 = 0;
    assign const_562_0 = 0;
    assign const_563_0 = 0;
    assign const_564_0 = 0;
    assign const_565_0 = 0;
    assign const_566_0 = 0;
    assign const_567_127 = 127;
    assign const_569_0 = 0;
    assign const_570_0 = 0;
    assign const_571_0 = 0;
    assign const_572_0 = 0;
    assign const_573_1 = 1;
    assign const_575_0 = 0;
    assign const_576_0 = 0;
    assign const_577_127 = 127;
    assign const_578_0 = 0;
    assign const_579_0 = 0;
    assign const_580_1 = 1;
    assign const_582_0 = 0;
    assign const_583_0 = 0;
    assign const_584_127 = 127;
    assign const_585_0 = 0;
    assign const_586_0 = 0;
    assign const_587_1 = 1;
    assign const_589_0 = 0;
    assign const_590_0 = 0;
    assign const_591_127 = 127;
    assign const_592_0 = 0;
    assign const_593_0 = 0;
    assign const_594_1 = 1;
    assign const_596_0 = 0;
    assign const_597_0 = 0;
    assign const_598_127 = 127;
    assign const_599_0 = 0;
    assign const_600_0 = 0;
    assign const_601_1 = 1;
    assign const_603_0 = 0;
    assign const_604_0 = 0;
    assign const_605_127 = 127;
    assign const_606_0 = 0;
    assign const_607_0 = 0;
    assign const_608_1 = 1;
    assign const_610_0 = 0;
    assign const_611_0 = 0;
    assign const_612_127 = 127;
    assign const_613_0 = 0;
    assign const_614_0 = 0;
    assign const_615_1 = 1;
    assign const_617_0 = 0;
    assign const_618_0 = 0;
    assign const_619_127 = 127;
    assign const_620_0 = 0;
    assign const_621_0 = 0;
    assign const_622_1 = 1;
    assign const_624_0 = 0;
    assign const_625_0 = 0;
    assign const_626_127 = 127;
    assign const_627_0 = 0;
    assign const_628_0 = 0;
    assign const_629_7 = 7;
    assign const_630_1 = 1;
    assign const_631_1 = 1;
    assign const_633_0 = 0;
    assign const_634_0 = 0;
    assign const_635_127 = 127;
    assign const_636_0 = 0;
    assign const_637_0 = 0;
    assign const_638_1 = 1;
    assign const_640_0 = 0;
    assign const_641_0 = 0;
    assign const_642_127 = 127;
    assign const_643_0 = 0;
    assign const_644_0 = 0;
    assign const_645_1 = 1;
    assign const_647_0 = 0;
    assign const_648_0 = 0;
    assign const_649_127 = 127;
    assign const_650_0 = 0;
    assign const_651_0 = 0;
    assign const_652_1 = 1;
    assign const_654_0 = 0;
    assign const_655_0 = 0;
    assign const_656_127 = 127;
    assign const_657_0 = 0;
    assign const_658_0 = 0;
    assign const_659_1 = 1;
    assign const_661_0 = 0;
    assign const_662_0 = 0;
    assign const_663_127 = 127;
    assign const_664_0 = 0;
    assign const_665_0 = 0;
    assign const_666_1 = 1;
    assign const_668_0 = 0;
    assign const_669_0 = 0;
    assign const_670_127 = 127;
    assign const_671_0 = 0;
    assign const_672_0 = 0;
    assign const_673_1 = 1;
    assign const_675_0 = 0;
    assign const_676_0 = 0;
    assign const_677_127 = 127;
    assign const_678_0 = 0;
    assign const_679_0 = 0;
    assign const_680_1 = 1;
    assign const_682_0 = 0;
    assign const_683_0 = 0;
    assign const_684_127 = 127;
    assign const_685_0 = 0;
    assign const_686_0 = 0;
    assign const_687_3 = 3;
    assign const_688_1 = 1;
    assign const_689_0 = 0;
    assign const_690_0 = 0;
    assign const_691_0 = 0;
    assign const_692_0 = 0;
    assign const_693_0 = 0;
    assign const_694_127 = 127;
    assign const_696_0 = 0;
    assign const_697_0 = 0;
    assign const_698_0 = 0;
    assign const_699_0 = 0;
    assign const_700_0 = 0;
    assign const_701_127 = 127;
    assign const_703_0 = 0;
    assign const_704_0 = 0;
    assign const_705_0 = 0;
    assign const_706_0 = 0;
    assign const_707_0 = 0;
    assign const_708_127 = 127;
    assign const_710_0 = 0;
    assign const_711_0 = 0;
    assign const_712_0 = 0;
    assign const_713_0 = 0;
    assign const_714_0 = 0;
    assign const_715_127 = 127;
    assign const_717_0 = 0;
    assign const_718_0 = 0;
    assign const_719_0 = 0;
    assign const_720_0 = 0;
    assign const_721_0 = 0;
    assign const_722_0 = 0;
    assign const_723_0 = 0;
    assign const_724_0 = 0;
    assign const_725_0 = 0;
    assign const_726_0 = 0;
    assign const_727_0 = 0;
    assign const_728_0 = 0;
    assign const_729_0 = 0;
    assign const_730_0 = 0;
    assign const_731_0 = 0;
    assign const_732_0 = 0;
    assign const_733_0 = 0;
    assign const_734_0 = 0;
    assign const_735_0 = 0;
    assign const_736_0 = 0;
    assign const_737_0 = 0;
    assign const_738_0 = 0;
    assign const_739_0 = 0;
    assign const_740_1 = 1;
    assign const_741_0 = 0;
    assign const_742_2 = 2;
    assign const_743_0 = 0;
    assign const_744_3 = 3;
    assign const_745_0 = 0;
    assign const_746_15 = 15;
    assign const_747_4 = 4;
    assign const_748_0 = 0;
    assign const_749_5 = 5;
    assign const_750_0 = 0;
    assign const_751_6 = 6;
    assign const_752_0 = 0;
    assign const_753_7 = 7;
    assign const_754_0 = 0;
    assign const_755_15 = 15;
    assign const_756_8 = 8;
    assign const_757_6 = 6;
    assign const_758_0 = 0;
    assign const_759_7 = 7;
    assign const_760_0 = 0;
    assign const_761_15 = 15;
    assign const_762_1 = 1;
    assign const_763_0 = 0;
    assign const_764_4 = 4;
    assign const_765_8 = 8;
    assign const_766_1 = 1;
    assign const_767_0 = 0;
    assign const_768_2 = 2;
    assign const_769_0 = 0;
    assign const_770_6 = 6;
    assign const_771_3 = 3;
    assign const_772_0 = 0;
    assign const_773_6 = 6;
    assign const_778_0 = 0;
    assign const_779_0 = 0;
    assign const_780_0 = 0;
    assign const_781_0 = 0;
    assign blue_o = tmp7940;
    assign green_o = tmp7929;
    assign red_o = tmp7912;
    assign tmp1 = {const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0};
    assign tmp2 = {tmp1, const_1_1};
    assign tmp3 = tmp0 + tmp2;
    assign tmp4 = {tmp3[26], tmp3[25], tmp3[24], tmp3[23], tmp3[22], tmp3[21], tmp3[20], tmp3[19], tmp3[18], tmp3[17], tmp3[16], tmp3[15], tmp3[14], tmp3[13], tmp3[12], tmp3[11], tmp3[10], tmp3[9], tmp3[8], tmp3[7], tmp3[6], tmp3[5], tmp3[4], tmp3[3], tmp3[2], tmp3[1], tmp3[0]};
    assign tmp8 = {tmp0[25]};
    assign tmp9 = tmp5 == tmp8;
    assign tmp10 = ~tmp9;
    assign tmp33 = ~tmp7;
    assign tmp35 = {tmp6211, const_3_0};
    assign tmp36 = my_calculator_ctrl == tmp35;
    assign tmp37 = my_calculator_ctrl == const_5_4;
    assign tmp61 = tmp4442 & tmp37;
    assign tmp75 = {tmp6211, const_15_1};
    assign tmp76 = my_calculator_ctrl == tmp75;
    assign tmp85 = my_calculator_in_x == tmp1117;
    assign tmp86 = my_calculator_in_x == const_19_15;
    assign tmp94 = tmp1093 & tmp196;
    assign tmp122 = tmp94 & tmp86;
    assign tmp125 = my_calculator_in_x == tmp1165;
    assign tmp128 = my_calculator_in_x == tmp7904;
    assign tmp129 = tmp125 | tmp128;
    assign tmp132 = my_calculator_in_x == tmp7908;
    assign tmp133 = tmp129 | tmp132;
    assign tmp146 = ~tmp520;
    assign tmp156 = tmp1194 ^ tmp1196;
    assign tmp160 = tmp1605 & tmp1200;
    assign tmp171 = ~tmp5229;
    assign tmp177 = tmp5532 - tmp1176;
    assign tmp178 = {tmp177[8]};
    assign tmp186 = tmp1225 | tmp1226;
    assign tmp187 = tmp2784 & tmp186;
    assign tmp196 = ~tmp85;
    assign tmp201 = {tmp12[6], tmp12[5], tmp12[4], tmp12[3], tmp12[2], tmp12[1], tmp12[0]};
    assign tmp202 = {tmp201, const_33_0};
    assign tmp214 = tmp1614 ^ tmp235;
    assign tmp219 = tmp202 - tmp5532;
    assign tmp220 = {tmp219[8]};
    assign tmp222 = ~tmp249;
    assign tmp223 = tmp220 ^ tmp222;
    assign tmp226 = tmp223 ^ tmp171;
    assign tmp227 = tmp214 & tmp226;
    assign tmp232 = tmp12 - tmp5532;
    assign tmp235 = ~tmp1615;
    assign tmp244 = tmp5532 - tmp202;
    assign tmp245 = {tmp244[8]};
    assign tmp248 = tmp245 ^ tmp171;
    assign tmp249 = {tmp202[7]};
    assign tmp251 = tmp248 ^ tmp222;
    assign tmp252 = tmp5532 == tmp202;
    assign tmp253 = tmp251 | tmp252;
    assign tmp254 = tmp701 & tmp253;
    assign tmp255 = tmp227 ? const_38_127 : tmp202;
    assign tmp256 = tmp254 ? _ver_out_tmp_31 : tmp255;
    assign tmp268 = {tmp15[6], tmp15[5], tmp15[4], tmp15[3], tmp15[2], tmp15[1], tmp15[0]};
    assign tmp287 = {tmp1331[8]};
    assign tmp290 = tmp287 ^ tmp1362;
    assign tmp299 = tmp15 - tmp5532;
    assign tmp312 = {tmp7358[8]};
    assign tmp320 = tmp1363 | tmp7366;
    assign tmp334 = tmp444 & tmp133;
    assign tmp345 = tmp897 ^ tmp171;
    assign tmp354 = {tmp7409[8]};
    assign tmp388 = tmp2320 & tmp7443;
    assign tmp404 = my_calculator_in_x == tmp1452;
    assign tmp407 = my_calculator_in_x == tmp1455;
    assign tmp408 = tmp404 | tmp407;
    assign tmp421 = tmp1099 & tmp408;
    assign tmp444 = tmp94 & tmp1046;
    assign tmp445 = ~tmp133;
    assign tmp514 = {const_59_0, const_58_4};
    assign tmp515 = my_calculator_in_x == tmp514;
    assign tmp518 = my_calculator_in_x == tmp7917;
    assign tmp519 = tmp515 | tmp518;
    assign tmp520 = {tmp11[7]};
    assign tmp526 = tmp1587 + tmp1712;
    assign tmp527 = {tmp526[8], tmp526[7], tmp526[6], tmp526[5], tmp526[4], tmp526[3], tmp526[2], tmp526[1], tmp526[0]};
    assign tmp528 = {tmp527[7], tmp527[6], tmp527[5], tmp527[4], tmp527[3], tmp527[2], tmp527[1], tmp527[0]};
    assign tmp549 = tmp1251 ^ tmp171;
    assign tmp550 = {tmp13[7]};
    assign tmp553 = tmp1605 & tmp1730;
    assign tmp558 = tmp528 - tmp5532;
    assign tmp559 = {tmp558[8]};
    assign tmp562 = tmp559 ^ tmp604;
    assign tmp565 = tmp562 ^ tmp171;
    assign tmp566 = tmp528 == tmp5532;
    assign tmp567 = tmp565 | tmp566;
    assign tmp568 = tmp553 & tmp567;
    assign tmp573 = tmp11 - tmp5532;
    assign tmp592 = tmp1279 ^ tmp171;
    assign tmp593 = tmp2784 & tmp592;
    assign tmp598 = tmp5532 - tmp528;
    assign tmp599 = {tmp598[8]};
    assign tmp602 = tmp599 ^ tmp171;
    assign tmp603 = {tmp528[7]};
    assign tmp604 = ~tmp603;
    assign tmp605 = tmp602 ^ tmp604;
    assign tmp607 = tmp605 | tmp566;
    assign tmp608 = tmp593 & tmp607;
    assign tmp609 = tmp568 ? const_68_127 : tmp528;
    assign tmp610 = tmp608 ? _ver_out_tmp_80 : tmp609;
    assign tmp644 = {tmp14[7]};
    assign tmp646 = {tmp644, tmp14};
    assign tmp647 = tmp1590 + tmp646;
    assign tmp648 = {tmp647[8], tmp647[7], tmp647[6], tmp647[5], tmp647[4], tmp647[3], tmp647[2], tmp647[1], tmp647[0]};
    assign tmp649 = {tmp648[7], tmp648[6], tmp648[5], tmp648[4], tmp648[3], tmp648[2], tmp648[1], tmp648[0]};
    assign tmp674 = tmp214 & tmp1742;
    assign tmp679 = tmp649 - tmp5532;
    assign tmp680 = {tmp679[8]};
    assign tmp681 = {tmp649[7]};
    assign tmp682 = ~tmp681;
    assign tmp683 = tmp680 ^ tmp682;
    assign tmp686 = tmp683 ^ tmp171;
    assign tmp687 = tmp649 == tmp5532;
    assign tmp688 = tmp686 | tmp687;
    assign tmp689 = tmp674 & tmp688;
    assign tmp698 = tmp2214 ^ tmp235;
    assign tmp701 = tmp698 ^ tmp171;
    assign tmp714 = tmp701 & tmp2271;
    assign tmp719 = tmp5532 - tmp649;
    assign tmp720 = {tmp719[8]};
    assign tmp723 = tmp720 ^ tmp171;
    assign tmp726 = tmp723 ^ tmp682;
    assign tmp728 = tmp726 | tmp687;
    assign tmp729 = tmp714 & tmp728;
    assign tmp730 = tmp689 ? const_76_127 : tmp649;
    assign tmp731 = tmp729 ? _ver_out_tmp_35 : tmp730;
    assign tmp768 = tmp1837 + tmp1962;
    assign tmp769 = {tmp768[8], tmp768[7], tmp768[6], tmp768[5], tmp768[4], tmp768[3], tmp768[2], tmp768[1], tmp768[0]};
    assign tmp770 = {tmp769[7], tmp769[6], tmp769[5], tmp769[4], tmp769[3], tmp769[2], tmp769[1], tmp769[0]};
    assign tmp795 = tmp1326 & tmp1980;
    assign tmp800 = tmp770 - tmp5532;
    assign tmp801 = {tmp800[8]};
    assign tmp803 = ~tmp845;
    assign tmp804 = tmp801 ^ tmp803;
    assign tmp807 = tmp804 ^ tmp171;
    assign tmp808 = tmp770 == tmp5532;
    assign tmp809 = tmp807 | tmp808;
    assign tmp810 = tmp795 & tmp809;
    assign tmp819 = tmp1889 ^ tmp7327;
    assign tmp835 = tmp2628 & tmp1420;
    assign tmp840 = tmp5532 - tmp770;
    assign tmp841 = {tmp840[8]};
    assign tmp844 = tmp841 ^ tmp171;
    assign tmp845 = {tmp770[7]};
    assign tmp847 = tmp844 ^ tmp803;
    assign tmp849 = tmp847 | tmp808;
    assign tmp850 = tmp835 & tmp849;
    assign tmp851 = tmp810 ? const_84_127 : tmp770;
    assign tmp852 = tmp850 ? _ver_out_tmp_38 : tmp851;
    assign tmp888 = {tmp7162, tmp18};
    assign tmp889 = tmp1840 + tmp888;
    assign tmp890 = {tmp889[8], tmp889[7], tmp889[6], tmp889[5], tmp889[4], tmp889[3], tmp889[2], tmp889[1], tmp889[0]};
    assign tmp891 = {tmp890[7], tmp890[6], tmp890[5], tmp890[4], tmp890[3], tmp890[2], tmp890[1], tmp890[0]};
    assign tmp897 = {tmp1860[8]};
    assign tmp902 = ~tmp938;
    assign tmp909 = {tmp6845[8]};
    assign tmp912 = tmp909 ^ tmp171;
    assign tmp916 = tmp7404 & tmp7556;
    assign tmp921 = tmp891 - tmp5532;
    assign tmp922 = {tmp921[8]};
    assign tmp923 = {tmp891[7]};
    assign tmp924 = ~tmp923;
    assign tmp925 = tmp922 ^ tmp924;
    assign tmp928 = tmp925 ^ tmp171;
    assign tmp930 = tmp928 | tmp969;
    assign tmp931 = tmp916 & tmp930;
    assign tmp937 = {tmp7422[8]};
    assign tmp938 = {tmp16[7]};
    assign tmp956 = tmp2320 & tmp2032;
    assign tmp961 = tmp5532 - tmp891;
    assign tmp962 = {tmp961[8]};
    assign tmp965 = tmp962 ^ tmp171;
    assign tmp968 = tmp965 ^ tmp924;
    assign tmp969 = tmp5532 == tmp891;
    assign tmp970 = tmp968 | tmp969;
    assign tmp971 = tmp956 & tmp970;
    assign tmp972 = tmp931 ? const_92_127 : tmp891;
    assign tmp973 = tmp971 ? _ver_out_tmp_40 : tmp972;
    assign tmp988 = tmp1101 & tmp519;
    assign tmp1004 = my_calculator_in_x == const_94_8;
    assign tmp1005 = tmp11 == _ver_out_tmp_41;
    assign tmp1028 = tmp1101 & tmp1077;
    assign tmp1030 = tmp12 == _ver_out_tmp_44;
    assign tmp1046 = ~tmp86;
    assign tmp1062 = {tmp6744[7], tmp6744[6], tmp6744[5], tmp6744[4], tmp6744[3], tmp6744[2], tmp6744[1], tmp6744[0]};
    assign tmp1077 = ~tmp519;
    assign tmp1093 = tmp3298 & tmp76;
    assign tmp1099 = tmp444 & tmp445;
    assign tmp1100 = ~tmp408;
    assign tmp1101 = tmp1099 & tmp1100;
    assign tmp1104 = tmp1028 & tmp1004;
    assign tmp1106 = {const_116_0, const_115_2};
    assign tmp1107 = my_calculator_ctrl == tmp1106;
    assign tmp1111 = ~tmp37;
    assign tmp1117 = {tmp1164, const_117_0};
    assign tmp1118 = my_calculator_in_y == tmp1117;
    assign tmp1119 = my_calculator_in_y == const_119_15;
    assign tmp1127 = tmp7644 & tmp1107;
    assign tmp1141 = tmp1240 & tmp1119;
    assign tmp1164 = {const_121_0, const_121_0, const_121_0};
    assign tmp1165 = {tmp1164, const_120_1};
    assign tmp1166 = my_calculator_in_y == tmp1165;
    assign tmp1169 = my_calculator_in_y == tmp7904;
    assign tmp1170 = tmp1166 | tmp1169;
    assign tmp1173 = my_calculator_in_y == tmp7908;
    assign tmp1174 = tmp1170 | tmp1173;
    assign tmp1175 = {tmp11[6], tmp11[5], tmp11[4], tmp11[3], tmp11[2], tmp11[1], tmp11[0]};
    assign tmp1176 = {tmp1175, const_126_0};
    assign tmp1181 = tmp5532 - tmp11;
    assign tmp1182 = {tmp1181[8]};
    assign tmp1193 = tmp1176 - tmp5532;
    assign tmp1194 = {tmp1193[8]};
    assign tmp1196 = ~tmp1223;
    assign tmp1200 = tmp156 ^ tmp171;
    assign tmp1222 = tmp178 ^ tmp171;
    assign tmp1223 = {tmp1176[7]};
    assign tmp1225 = tmp1222 ^ tmp1196;
    assign tmp1226 = tmp5532 == tmp1176;
    assign tmp1229 = tmp160 ? const_131_127 : tmp1176;
    assign tmp1230 = tmp187 ? _ver_out_tmp_28 : tmp1229;
    assign tmp1240 = tmp1127 & tmp1496;
    assign tmp1244 = {tmp13[6], tmp13[5], tmp13[4], tmp13[3], tmp13[2], tmp13[1], tmp13[0]};
    assign tmp1245 = {tmp1244, const_133_0};
    assign tmp1250 = tmp5532 - tmp13;
    assign tmp1251 = {tmp1250[8]};
    assign tmp1262 = tmp1245 - tmp5532;
    assign tmp1263 = {tmp1262[8]};
    assign tmp1264 = {tmp1245[7]};
    assign tmp1266 = tmp1263 ^ tmp1293;
    assign tmp1269 = tmp1266 ^ tmp171;
    assign tmp1270 = tmp1730 & tmp1269;
    assign tmp1279 = tmp1764 ^ tmp2255;
    assign tmp1287 = tmp5532 - tmp1245;
    assign tmp1288 = {tmp1287[8]};
    assign tmp1291 = tmp1288 ^ tmp171;
    assign tmp1293 = ~tmp1264;
    assign tmp1294 = tmp1291 ^ tmp1293;
    assign tmp1295 = tmp5532 == tmp1245;
    assign tmp1296 = tmp1294 | tmp1295;
    assign tmp1297 = tmp592 & tmp1296;
    assign tmp1298 = tmp1270 ? const_138_127 : tmp1245;
    assign tmp1299 = tmp1297 ? _ver_out_tmp_58 : tmp1298;
    assign tmp1320 = {tmp7321[8]};
    assign tmp1326 = tmp7325 ^ tmp7327;
    assign tmp1331 = tmp7316 - tmp5532;
    assign tmp1338 = tmp290 ^ tmp171;
    assign tmp1361 = {tmp7316[7]};
    assign tmp1362 = ~tmp1361;
    assign tmp1363 = tmp7362 ^ tmp1362;
    assign tmp1367 = tmp7341 ? const_145_127 : tmp7316;
    assign tmp1381 = tmp2159 & tmp1174;
    assign tmp1392 = tmp7474 ^ tmp171;
    assign tmp1400 = tmp7468 - tmp5532;
    assign tmp1404 = tmp7486 ^ tmp7488;
    assign tmp1407 = tmp1404 ^ tmp171;
    assign tmp1413 = tmp17 - tmp5532;
    assign tmp1420 = tmp7502 ^ tmp171;
    assign tmp1425 = tmp5532 - tmp7468;
    assign tmp1426 = {tmp1425[8]};
    assign tmp1429 = tmp1426 ^ tmp171;
    assign tmp1434 = tmp7517 | tmp7518;
    assign tmp1435 = tmp1420 & tmp1434;
    assign tmp1436 = tmp7493 ? const_152_127 : tmp7468;
    assign tmp1437 = tmp1435 ? _ver_out_tmp_63 : tmp1436;
    assign tmp1452 = {const_155_0, const_154_6};
    assign tmp1453 = my_calculator_in_y == tmp1452;
    assign tmp1455 = {const_157_0, const_156_7};
    assign tmp1456 = my_calculator_in_y == tmp1455;
    assign tmp1457 = tmp1453 | tmp1456;
    assign tmp1468 = ~tmp1119;
    assign tmp1496 = ~tmp1118;
    assign tmp1548 = ~tmp33;
    assign tmp1577 = tmp2188 & tmp1457;
    assign tmp1580 = my_calculator_in_y == tmp514;
    assign tmp1583 = my_calculator_in_y == tmp7917;
    assign tmp1584 = tmp1580 | tmp1583;
    assign tmp1587 = {tmp520, tmp11};
    assign tmp1590 = {tmp1615, tmp12};
    assign tmp1591 = tmp1587 + tmp1590;
    assign tmp1592 = {tmp1591[8], tmp1591[7], tmp1591[6], tmp1591[5], tmp1591[4], tmp1591[3], tmp1591[2], tmp1591[1], tmp1591[0]};
    assign tmp1593 = {tmp1592[7], tmp1592[6], tmp1592[5], tmp1592[4], tmp1592[3], tmp1592[2], tmp1592[1], tmp1592[0]};
    assign tmp1602 = tmp1182 ^ tmp171;
    assign tmp1605 = tmp1602 ^ tmp146;
    assign tmp1611 = {tmp6763[8]};
    assign tmp1614 = tmp1611 ^ tmp171;
    assign tmp1615 = {tmp12[7]};
    assign tmp1618 = tmp1605 & tmp214;
    assign tmp1623 = tmp1593 - tmp5532;
    assign tmp1624 = {tmp1623[8]};
    assign tmp1625 = {tmp1593[7]};
    assign tmp1626 = ~tmp1625;
    assign tmp1627 = tmp1624 ^ tmp1626;
    assign tmp1630 = tmp1627 ^ tmp171;
    assign tmp1632 = tmp1630 | tmp1671;
    assign tmp1633 = tmp1618 & tmp1632;
    assign tmp1658 = tmp2784 & tmp701;
    assign tmp1663 = tmp5532 - tmp1593;
    assign tmp1664 = {tmp1663[8]};
    assign tmp1667 = tmp1664 ^ tmp171;
    assign tmp1670 = tmp1667 ^ tmp1626;
    assign tmp1671 = tmp5532 == tmp1593;
    assign tmp1672 = tmp1670 | tmp1671;
    assign tmp1673 = tmp1658 & tmp1672;
    assign tmp1674 = tmp1633 ? const_168_127 : tmp1593;
    assign tmp1675 = tmp1673 ? _ver_out_tmp_67 : tmp1674;
    assign tmp1709 = tmp2190 & tmp1584;
    assign tmp1712 = {tmp550, tmp13};
    assign tmp1716 = tmp1712 + tmp646;
    assign tmp1717 = {tmp1716[8], tmp1716[7], tmp1716[6], tmp1716[5], tmp1716[4], tmp1716[3], tmp1716[2], tmp1716[1], tmp1716[0]};
    assign tmp1718 = {tmp1717[7], tmp1717[6], tmp1717[5], tmp1717[4], tmp1717[3], tmp1717[2], tmp1717[1], tmp1717[0]};
    assign tmp1730 = tmp549 ^ tmp2255;
    assign tmp1735 = tmp5532 - tmp14;
    assign tmp1736 = {tmp1735[8]};
    assign tmp1739 = tmp1736 ^ tmp171;
    assign tmp1742 = tmp1739 ^ tmp1778;
    assign tmp1743 = tmp1730 & tmp1742;
    assign tmp1748 = tmp1718 - tmp5532;
    assign tmp1749 = {tmp1748[8]};
    assign tmp1750 = {tmp1718[7]};
    assign tmp1752 = tmp1749 ^ tmp1794;
    assign tmp1755 = tmp1752 ^ tmp171;
    assign tmp1756 = tmp1718 == tmp5532;
    assign tmp1757 = tmp1755 | tmp1756;
    assign tmp1758 = tmp1743 & tmp1757;
    assign tmp1763 = tmp13 - tmp5532;
    assign tmp1764 = {tmp1763[8]};
    assign tmp1776 = {tmp2264[8]};
    assign tmp1778 = ~tmp644;
    assign tmp1783 = tmp592 & tmp2271;
    assign tmp1788 = tmp5532 - tmp1718;
    assign tmp1789 = {tmp1788[8]};
    assign tmp1792 = tmp1789 ^ tmp171;
    assign tmp1794 = ~tmp1750;
    assign tmp1795 = tmp1792 ^ tmp1794;
    assign tmp1797 = tmp1795 | tmp1756;
    assign tmp1798 = tmp1783 & tmp1797;
    assign tmp1799 = tmp1758 ? const_176_127 : tmp1718;
    assign tmp1800 = tmp1798 ? _ver_out_tmp_10 : tmp1799;
    assign tmp1815 = ~tmp1457;
    assign tmp1837 = {tmp2623, tmp15};
    assign tmp1840 = {tmp938, tmp16};
    assign tmp1841 = tmp1837 + tmp1840;
    assign tmp1842 = {tmp1841[8], tmp1841[7], tmp1841[6], tmp1841[5], tmp1841[4], tmp1841[3], tmp1841[2], tmp1841[1], tmp1841[0]};
    assign tmp1843 = {tmp1842[7], tmp1842[6], tmp1842[5], tmp1842[4], tmp1842[3], tmp1842[2], tmp1842[1], tmp1842[0]};
    assign tmp1860 = tmp5532 - tmp16;
    assign tmp1868 = tmp1326 & tmp7404;
    assign tmp1873 = tmp1843 - tmp5532;
    assign tmp1874 = {tmp1873[8]};
    assign tmp1876 = ~tmp1918;
    assign tmp1877 = tmp1874 ^ tmp1876;
    assign tmp1880 = tmp1877 ^ tmp171;
    assign tmp1882 = tmp1880 | tmp1921;
    assign tmp1883 = tmp1868 & tmp1882;
    assign tmp1889 = {tmp299[8]};
    assign tmp1904 = tmp937 ^ tmp902;
    assign tmp1908 = tmp2628 & tmp2320;
    assign tmp1913 = tmp5532 - tmp1843;
    assign tmp1914 = {tmp1913[8]};
    assign tmp1917 = tmp1914 ^ tmp171;
    assign tmp1918 = {tmp1843[7]};
    assign tmp1920 = tmp1917 ^ tmp1876;
    assign tmp1921 = tmp5532 == tmp1843;
    assign tmp1922 = tmp1920 | tmp1921;
    assign tmp1923 = tmp1908 & tmp1922;
    assign tmp1924 = tmp1883 ? const_184_127 : tmp1843;
    assign tmp1925 = tmp1923 ? _ver_out_tmp_71 : tmp1924;
    assign tmp1962 = {tmp7121, tmp17};
    assign tmp1966 = tmp1962 + tmp888;
    assign tmp1967 = {tmp1966[8], tmp1966[7], tmp1966[6], tmp1966[5], tmp1966[4], tmp1966[3], tmp1966[2], tmp1966[1], tmp1966[0]};
    assign tmp1968 = {tmp1967[7], tmp1967[6], tmp1967[5], tmp1967[4], tmp1967[3], tmp1967[2], tmp1967[1], tmp1967[0]};
    assign tmp1973 = tmp5532 - tmp17;
    assign tmp1979 = ~tmp7121;
    assign tmp1980 = tmp1392 ^ tmp1979;
    assign tmp1993 = tmp1980 & tmp7556;
    assign tmp1998 = tmp1968 - tmp5532;
    assign tmp1999 = {tmp1998[8]};
    assign tmp2000 = {tmp1968[7]};
    assign tmp2001 = ~tmp2000;
    assign tmp2002 = tmp1999 ^ tmp2001;
    assign tmp2005 = tmp2002 ^ tmp171;
    assign tmp2007 = tmp2005 | tmp2046;
    assign tmp2008 = tmp1993 & tmp2007;
    assign tmp2014 = {tmp1413[8]};
    assign tmp2026 = {tmp2351[8]};
    assign tmp2032 = tmp2355 ^ tmp171;
    assign tmp2033 = tmp1420 & tmp2032;
    assign tmp2038 = tmp5532 - tmp1968;
    assign tmp2039 = {tmp2038[8]};
    assign tmp2042 = tmp2039 ^ tmp171;
    assign tmp2045 = tmp2042 ^ tmp2001;
    assign tmp2046 = tmp5532 == tmp1968;
    assign tmp2047 = tmp2045 | tmp2046;
    assign tmp2048 = tmp2033 & tmp2047;
    assign tmp2049 = tmp2008 ? const_192_127 : tmp1968;
    assign tmp2050 = tmp2048 ? _ver_out_tmp_73 : tmp2049;
    assign tmp2085 = my_calculator_in_y == const_194_8;
    assign tmp2095 = ~tmp36;
    assign tmp2113 = tmp13 == _ver_out_tmp_77;
    assign tmp2120 = {tmp2877[7], tmp2877[6], tmp2877[5], tmp2877[4], tmp2877[3], tmp2877[2], tmp2877[1], tmp2877[0]};
    assign tmp2138 = tmp2190 & tmp2164;
    assign tmp2159 = tmp1240 & tmp1468;
    assign tmp2164 = ~tmp1584;
    assign tmp2174 = {tmp6813[7], tmp6813[6], tmp6813[5], tmp6813[4], tmp6813[3], tmp6813[2], tmp6813[1], tmp6813[0]};
    assign tmp2187 = ~tmp1174;
    assign tmp2188 = tmp2159 & tmp2187;
    assign tmp2190 = tmp2188 & tmp1815;
    assign tmp2193 = tmp2138 & tmp2085;
    assign tmp2195 = {const_216_0, const_215_3};
    assign tmp2196 = my_calculator_ctrl == tmp2195;
    assign tmp2214 = {tmp232[8]};
    assign tmp2221 = tmp2784 == tmp701;
    assign tmp2246 = tmp701 == tmp592;
    assign tmp2247 = tmp2221 & tmp2246;
    assign tmp2255 = ~tmp550;
    assign tmp2264 = tmp14 - tmp5532;
    assign tmp2268 = tmp1776 ^ tmp1778;
    assign tmp2271 = tmp2268 ^ tmp171;
    assign tmp2272 = tmp592 == tmp2271;
    assign tmp2273 = tmp2247 & tmp2272;
    assign tmp2308 = tmp2628 == tmp2320;
    assign tmp2320 = tmp1904 ^ tmp171;
    assign tmp2333 = tmp2320 == tmp1420;
    assign tmp2334 = tmp2308 & tmp2333;
    assign tmp2351 = tmp18 - tmp5532;
    assign tmp2354 = ~tmp7162;
    assign tmp2355 = tmp2026 ^ tmp2354;
    assign tmp2359 = tmp1420 == tmp2032;
    assign tmp2360 = tmp2334 & tmp2359;
    assign tmp2377 = tmp2738 | tmp2741;
    assign tmp2380 = tmp17 == tmp5532;
    assign tmp2381 = tmp2377 | tmp2380;
    assign tmp2384 = tmp18 == tmp5532;
    assign tmp2385 = tmp2381 | tmp2384;
    assign tmp2396 = tmp7845 & tmp7846;
    assign tmp2397 = ~tmp7847;
    assign tmp2398 = tmp2396 & tmp2397;
    assign tmp2409 = {tmp11[0]};
    assign tmp2410 = {tmp12[0]};
    assign tmp2411 = tmp2409 | tmp2410;
    assign tmp2412 = {tmp13[0]};
    assign tmp2413 = tmp2411 | tmp2412;
    assign tmp2414 = {tmp14[0]};
    assign tmp2415 = tmp2413 | tmp2414;
    assign tmp2416 = ~tmp2415;
    assign tmp2432 = {tmp573[8]};
    assign tmp2439 = tmp7848 & tmp2784;
    assign tmp2452 = tmp2439 & tmp2628;
    assign tmp2459 = tmp1005 ? tmp2534 : tmp1181;
    assign tmp2460 = {tmp2459[7], tmp2459[6], tmp2459[5], tmp2459[4], tmp2459[3], tmp2459[2], tmp2459[1], tmp2459[0]};
    assign tmp2516 = tmp6830 ? tmp2534 : tmp1735;
    assign tmp2517 = {tmp2516[7], tmp2516[6], tmp2516[5], tmp2516[4], tmp2516[3], tmp2516[2], tmp2516[1], tmp2516[0]};
    assign tmp2534 = {tmp6211, const_262_127};
    assign tmp2548 = tmp16 == _ver_out_tmp_5;
    assign tmp2555 = {tmp7088[7], tmp7088[6], tmp7088[5], tmp7088[4], tmp7088[3], tmp7088[2], tmp7088[1], tmp7088[0]};
    assign tmp2566 = tmp2706 & tmp2452;
    assign tmp2586 = tmp18 == _ver_out_tmp_8;
    assign tmp2593 = {tmp6848[7], tmp6848[6], tmp6848[5], tmp6848[4], tmp6848[3], tmp6848[2], tmp6848[1], tmp6848[0]};
    assign tmp2623 = {tmp15[7]};
    assign tmp2628 = tmp819 ^ tmp171;
    assign tmp2629 = tmp2784 & tmp2628;
    assign tmp2630 = ~tmp2629;
    assign tmp2631 = tmp7848 & tmp2630;
    assign tmp2702 = ~tmp76;
    assign tmp2706 = tmp3157 & tmp2196;
    assign tmp2730 = ~tmp1107;
    assign tmp2733 = ~tmp2452;
    assign tmp2734 = tmp2706 & tmp2733;
    assign tmp2735 = tmp2734 & tmp2631;
    assign tmp2736 = {const_282_0, const_282_0, const_282_0, const_282_0, const_282_0, const_282_0, const_282_0};
    assign tmp2738 = tmp15 == tmp5532;
    assign tmp2741 = tmp16 == tmp5532;
    assign tmp2742 = tmp2738 & tmp2741;
    assign tmp2746 = tmp2742 & tmp2380;
    assign tmp2750 = tmp2746 & tmp2384;
    assign tmp2772 = tmp2706 & tmp2750;
    assign tmp2781 = tmp2432 ^ tmp146;
    assign tmp2784 = tmp2781 ^ tmp171;
    assign tmp2797 = tmp2784 == tmp2628;
    assign tmp2798 = ~tmp2797;
    assign tmp2856 = {tmp6766[7], tmp6766[6], tmp6766[5], tmp6766[4], tmp6766[3], tmp6766[2], tmp6766[1], tmp6766[0]};
    assign tmp2877 = tmp2113 ? tmp2534 : tmp1250;
    assign tmp2892 = tmp5355 & tmp2798;
    assign tmp2916 = {tmp4817[6]};
    assign tmp2921 = tmp7869 - tmp3588;
    assign tmp2922 = {tmp2921[8]};
    assign tmp2923 = {tmp3588[7]};
    assign tmp2924 = ~tmp2923;
    assign tmp2925 = tmp2922 ^ tmp2924;
    assign tmp2928 = tmp2925 ^ tmp5510;
    assign tmp2929 = tmp3588 == tmp7869;
    assign tmp2930 = tmp2928 | tmp2929;
    assign tmp2937 = tmp7873 - tmp3038;
    assign tmp2938 = {tmp2937[8]};
    assign tmp2941 = tmp2938 ^ tmp3609;
    assign tmp2944 = tmp2941 ^ tmp3554;
    assign tmp2945 = tmp3038 == tmp7873;
    assign tmp2946 = tmp2944 | tmp2945;
    assign tmp2947 = tmp2930 & tmp2946;
    assign tmp2948 = {tmp7861[7], tmp7861[6], tmp7861[5], tmp7861[4], tmp7861[3], tmp7861[2], tmp7861[1]};
    assign tmp2954 = tmp7877 - tmp4876;
    assign tmp2955 = {tmp2954[8]};
    assign tmp2958 = tmp2955 ^ tmp3624;
    assign tmp2961 = tmp2958 ^ tmp4246;
    assign tmp2962 = tmp4876 == tmp7877;
    assign tmp2963 = tmp2961 | tmp2962;
    assign tmp2964 = tmp2947 & tmp2963;
    assign tmp2971 = tmp7881 - tmp3633;
    assign tmp2972 = {tmp2971[8]};
    assign tmp2974 = ~tmp3638;
    assign tmp2975 = tmp2972 ^ tmp2974;
    assign tmp2978 = tmp2975 ^ tmp4698;
    assign tmp2979 = tmp3633 == tmp7881;
    assign tmp2980 = tmp2978 | tmp2979;
    assign tmp2981 = tmp2964 & tmp2980;
    assign tmp3036 = {tmp4845[6]};
    assign tmp3038 = {tmp3036, tmp4845};
    assign tmp3055 = tmp3113 & tmp7849;
    assign tmp3077 = {tmp7865[7], tmp7865[6], tmp7865[5], tmp7865[4], tmp7865[3], tmp7865[2], tmp7865[1]};
    assign tmp3078 = {tmp3077[6]};
    assign tmp3113 = tmp4274 & tmp2981;
    assign tmp3157 = tmp7644 & tmp2730;
    assign tmp3194 = ~tmp2750;
    assign tmp3197 = ~tmp2798;
    assign tmp3201 = tmp3113 & tmp5447;
    assign tmp3238 = {tmp7869[6], tmp7869[5], tmp7869[4], tmp7869[3], tmp7869[2], tmp7869[1], tmp7869[0]};
    assign tmp3239 = {tmp3238, const_317_0};
    assign tmp3245 = {tmp5521[8]};
    assign tmp3260 = tmp5144 ^ tmp5146;
    assign tmp3270 = {tmp5546[8]};
    assign tmp3282 = {tmp5168[8]};
    assign tmp3285 = tmp3282 ^ tmp171;
    assign tmp3286 = {tmp3239[7]};
    assign tmp3288 = tmp3285 ^ tmp5146;
    assign tmp3290 = tmp3288 | tmp5176;
    assign tmp3291 = tmp5553 & tmp3290;
    assign tmp3298 = tmp4442 & tmp1111;
    assign tmp3319 = {tmp6210[8]};
    assign tmp3322 = tmp3319 ^ tmp171;
    assign tmp3350 = tmp4583 ^ tmp171;
    assign tmp3366 = tmp5232 ? const_329_127 : tmp5207;
    assign tmp3367 = tmp5259 ? _ver_out_tmp_29 : tmp3366;
    assign tmp3404 = tmp5784 - tmp5532;
    assign tmp3417 = tmp7877 - tmp5532;
    assign tmp3421 = tmp5815 ^ tmp4246;
    assign tmp3429 = tmp5532 - tmp5784;
    assign tmp3430 = {tmp3429[8]};
    assign tmp3433 = tmp3430 ^ tmp171;
    assign tmp3435 = ~tmp5831;
    assign tmp3436 = tmp3433 ^ tmp3435;
    assign tmp3438 = tmp3436 | tmp5834;
    assign tmp3440 = tmp5313 ? const_336_127 : tmp5784;
    assign tmp3460 = {tmp7881[6], tmp7881[5], tmp7881[4], tmp7881[3], tmp7881[2], tmp7881[1], tmp7881[0]};
    assign tmp3461 = {tmp3460, const_338_0};
    assign tmp3470 = tmp4711 ^ tmp171;
    assign tmp3473 = tmp3470 ^ tmp4698;
    assign tmp3486 = tmp3473 & tmp5942;
    assign tmp3491 = tmp7881 - tmp5532;
    assign tmp3492 = {tmp3491[8]};
    assign tmp3495 = tmp3492 ^ tmp4698;
    assign tmp3498 = tmp3495 ^ tmp171;
    assign tmp3504 = {tmp5960[8]};
    assign tmp3507 = tmp3504 ^ tmp171;
    assign tmp3511 = tmp5532 == tmp3461;
    assign tmp3512 = tmp5418 | tmp3511;
    assign tmp3515 = tmp5970 ? _ver_out_tmp_83 : tmp5971;
    assign tmp3537 = {tmp4462[8]};
    assign tmp3540 = tmp3537 ^ tmp3762;
    assign tmp3543 = tmp3540 ^ tmp5510;
    assign tmp3544 = tmp7853 == tmp7869;
    assign tmp3545 = tmp3543 | tmp3544;
    assign tmp3551 = ~tmp3895;
    assign tmp3552 = tmp4540 ^ tmp3551;
    assign tmp3554 = ~tmp5660;
    assign tmp3555 = tmp3552 ^ tmp3554;
    assign tmp3556 = tmp7857 == tmp7873;
    assign tmp3557 = tmp3555 | tmp3556;
    assign tmp3558 = tmp3545 & tmp3557;
    assign tmp3562 = {tmp4617[8]};
    assign tmp3565 = tmp3562 ^ tmp4623;
    assign tmp3568 = tmp3565 ^ tmp4246;
    assign tmp3569 = tmp7861 == tmp7877;
    assign tmp3570 = tmp3568 | tmp3569;
    assign tmp3571 = tmp3558 & tmp3570;
    assign tmp3574 = tmp7881 - tmp7865;
    assign tmp3575 = {tmp3574[8]};
    assign tmp3578 = tmp3575 ^ tmp4164;
    assign tmp3579 = {tmp7881[7]};
    assign tmp3581 = tmp3578 ^ tmp4698;
    assign tmp3582 = tmp7865 == tmp7881;
    assign tmp3583 = tmp3581 | tmp3582;
    assign tmp3584 = tmp3571 & tmp3583;
    assign tmp3588 = {tmp2916, tmp4817};
    assign tmp3591 = tmp3588 - tmp7869;
    assign tmp3592 = {tmp3591[8]};
    assign tmp3595 = tmp3592 ^ tmp2924;
    assign tmp3598 = tmp3595 ^ tmp5510;
    assign tmp3599 = tmp3584 & tmp3598;
    assign tmp3606 = tmp3038 - tmp7873;
    assign tmp3607 = {tmp3606[8]};
    assign tmp3608 = {tmp3038[7]};
    assign tmp3609 = ~tmp3608;
    assign tmp3610 = tmp3607 ^ tmp3609;
    assign tmp3613 = tmp3610 ^ tmp3554;
    assign tmp3614 = tmp3599 & tmp3613;
    assign tmp3621 = tmp4876 - tmp7877;
    assign tmp3622 = {tmp3621[8]};
    assign tmp3623 = {tmp4876[7]};
    assign tmp3624 = ~tmp3623;
    assign tmp3625 = tmp3622 ^ tmp3624;
    assign tmp3628 = tmp3625 ^ tmp4246;
    assign tmp3629 = tmp3614 & tmp3628;
    assign tmp3633 = {tmp3078, tmp3077};
    assign tmp3636 = tmp3633 - tmp7881;
    assign tmp3637 = {tmp3636[8]};
    assign tmp3638 = {tmp3633[7]};
    assign tmp3640 = tmp3637 ^ tmp2974;
    assign tmp3643 = tmp3640 ^ tmp4698;
    assign tmp3644 = tmp3629 & tmp3643;
    assign tmp3698 = tmp4456 & tmp3644;
    assign tmp3699 = _ver_out_tmp_37 == tmp7869;
    assign tmp3705 = tmp3699 ? tmp2534 : tmp5521;
    assign tmp3708 = {tmp6067, tmp7853};
    assign tmp3711 = {tmp3736, tmp3705};
    assign tmp3712 = tmp3708 + tmp3711;
    assign tmp3713 = {tmp3712[9], tmp3712[8], tmp3712[7], tmp3712[6], tmp3712[5], tmp3712[4], tmp3712[3], tmp3712[2], tmp3712[1], tmp3712[0]};
    assign tmp3731 = tmp6533 - tmp3705;
    assign tmp3732 = {tmp3731[9]};
    assign tmp3735 = tmp3732 ^ tmp6538;
    assign tmp3736 = {tmp3705[8]};
    assign tmp3737 = ~tmp3736;
    assign tmp3738 = tmp3735 ^ tmp3737;
    assign tmp3739 = tmp5462 & tmp3738;
    assign tmp3746 = {tmp6074[7]};
    assign tmp3747 = ~tmp3746;
    assign tmp3748 = tmp6105 ^ tmp3747;
    assign tmp3752 = tmp6074 == tmp5532;
    assign tmp3753 = tmp6111 | tmp3752;
    assign tmp3754 = tmp3739 & tmp3753;
    assign tmp3759 = tmp7853 - tmp5532;
    assign tmp3760 = {tmp3759[8]};
    assign tmp3762 = ~tmp6084;
    assign tmp3771 = tmp3705 - tmp6533;
    assign tmp3775 = tmp6132 ^ tmp3737;
    assign tmp3794 = tmp6139 & tmp6153;
    assign tmp3795 = tmp3754 ? const_358_127 : tmp6074;
    assign tmp3833 = _ver_out_tmp_43 == tmp7873;
    assign tmp3841 = {tmp3895, tmp3895};
    assign tmp3842 = {tmp3841, tmp7857};
    assign tmp3845 = {tmp6244, tmp6213};
    assign tmp3846 = tmp3842 + tmp3845;
    assign tmp3853 = tmp5532 - tmp7857;
    assign tmp3854 = {tmp3853[8]};
    assign tmp3857 = tmp3854 ^ tmp171;
    assign tmp3865 = tmp6533 - tmp6213;
    assign tmp3878 = tmp6222 - tmp5532;
    assign tmp3893 = tmp7857 - tmp5532;
    assign tmp3894 = {tmp3893[8]};
    assign tmp3895 = {tmp7857[7]};
    assign tmp3897 = tmp3894 ^ tmp3551;
    assign tmp3906 = {tmp6279[9]};
    assign tmp3925 = tmp6296 ^ tmp6298;
    assign tmp3927 = tmp3925 | tmp6300;
    assign tmp3928 = tmp6287 & tmp3927;
    assign tmp3970 = tmp5532 - tmp7877;
    assign tmp3973 = tmp6355 ? tmp2534 : tmp3970;
    assign tmp3975 = {tmp5749, tmp5749};
    assign tmp3976 = {tmp3975, tmp7861};
    assign tmp3979 = {tmp4041, tmp3973};
    assign tmp3994 = tmp5726 ^ tmp4623;
    assign tmp3999 = tmp6533 - tmp3973;
    assign tmp4003 = tmp6388 ^ tmp6538;
    assign tmp4005 = ~tmp4041;
    assign tmp4007 = tmp3994 & tmp6394;
    assign tmp4021 = tmp6407 | tmp4060;
    assign tmp4040 = {tmp6427[9]};
    assign tmp4041 = {tmp3973[8]};
    assign tmp4043 = tmp4040 ^ tmp4005;
    assign tmp4046 = tmp4043 ^ tmp6538;
    assign tmp4047 = tmp6422 & tmp4046;
    assign tmp4053 = {tmp6440[8]};
    assign tmp4060 = tmp5532 == tmp6370;
    assign tmp4064 = tmp6450 ? _ver_out_tmp_1 : tmp6451;
    assign tmp4101 = _ver_out_tmp_2 == tmp7881;
    assign tmp4113 = {tmp6577, tmp6509};
    assign tmp4116 = {tmp6517[7], tmp6517[6], tmp6517[5], tmp6517[4], tmp6517[3], tmp6517[2], tmp6517[1], tmp6517[0]};
    assign tmp4121 = tmp5532 - tmp7865;
    assign tmp4122 = {tmp4121[8]};
    assign tmp4125 = tmp4122 ^ tmp171;
    assign tmp4134 = {tmp6535[9]};
    assign tmp4146 = tmp4116 - tmp5532;
    assign tmp4147 = {tmp4146[8]};
    assign tmp4149 = ~tmp4191;
    assign tmp4163 = {tmp7865[7]};
    assign tmp4164 = ~tmp4163;
    assign tmp4174 = {tmp6575[9]};
    assign tmp4180 = tmp6579 ^ tmp6538;
    assign tmp4187 = {tmp6588[8]};
    assign tmp4191 = {tmp4116[7]};
    assign tmp4194 = tmp5532 == tmp4116;
    assign tmp4198 = tmp6598 ? _ver_out_tmp_7 : tmp6599;
    assign tmp4219 = tmp7853 - tmp7869;
    assign tmp4220 = {tmp4219[8]};
    assign tmp4223 = tmp4220 ^ tmp3762;
    assign tmp4226 = tmp4223 ^ tmp5510;
    assign tmp4229 = tmp7857 - tmp7873;
    assign tmp4230 = {tmp4229[8]};
    assign tmp4233 = tmp4230 ^ tmp3551;
    assign tmp4236 = tmp4233 ^ tmp3554;
    assign tmp4237 = tmp4226 & tmp4236;
    assign tmp4240 = tmp7861 - tmp7877;
    assign tmp4241 = {tmp4240[8]};
    assign tmp4244 = tmp4241 ^ tmp4623;
    assign tmp4246 = ~tmp4619;
    assign tmp4247 = tmp4244 ^ tmp4246;
    assign tmp4248 = tmp4237 & tmp4247;
    assign tmp4251 = tmp7865 - tmp7881;
    assign tmp4252 = {tmp4251[8]};
    assign tmp4255 = tmp4252 ^ tmp4164;
    assign tmp4258 = tmp4255 ^ tmp4698;
    assign tmp4259 = tmp4248 & tmp4258;
    assign tmp4274 = tmp5355 & tmp3197;
    assign tmp4311 = tmp2706 & tmp3194;
    assign tmp4359 = tmp6670 & tmp4259;
    assign tmp4442 = tmp1548 & tmp2095;
    assign tmp4456 = tmp4274 & tmp4992;
    assign tmp4462 = tmp7869 - tmp7853;
    assign tmp4466 = tmp3537 ^ tmp5510;
    assign tmp4469 = tmp4466 ^ tmp3762;
    assign tmp4470 = {tmp7869[5], tmp7869[4], tmp7869[3], tmp7869[2], tmp7869[1], tmp7869[0]};
    assign tmp4471 = {tmp4470, const_401_0};
    assign tmp4488 = tmp4471 - tmp5532;
    assign tmp4489 = {tmp4488[8]};
    assign tmp4490 = {tmp4471[7]};
    assign tmp4492 = tmp4489 ^ tmp4519;
    assign tmp4495 = tmp4492 ^ tmp171;
    assign tmp4496 = tmp5528 & tmp4495;
    assign tmp4513 = tmp5532 - tmp4471;
    assign tmp4514 = {tmp4513[8]};
    assign tmp4517 = tmp4514 ^ tmp171;
    assign tmp4519 = ~tmp4490;
    assign tmp4520 = tmp4517 ^ tmp4519;
    assign tmp4521 = tmp5532 == tmp4471;
    assign tmp4522 = tmp4520 | tmp4521;
    assign tmp4523 = tmp5553 & tmp4522;
    assign tmp4524 = tmp4496 ? const_406_127 : tmp4471;
    assign tmp4525 = tmp4523 ? _ver_out_tmp_9 : tmp4524;
    assign tmp4528 = tmp7853 - tmp4525;
    assign tmp4529 = {tmp4528[8]};
    assign tmp4532 = tmp4529 ^ tmp3762;
    assign tmp4533 = {tmp4525[7]};
    assign tmp4534 = ~tmp4533;
    assign tmp4535 = tmp4532 ^ tmp4534;
    assign tmp4536 = tmp4469 & tmp4535;
    assign tmp4539 = tmp7873 - tmp7857;
    assign tmp4540 = {tmp4539[8]};
    assign tmp4543 = tmp4540 ^ tmp3554;
    assign tmp4546 = tmp4543 ^ tmp3551;
    assign tmp4547 = tmp4536 & tmp4546;
    assign tmp4548 = {tmp7873[5], tmp7873[4], tmp7873[3], tmp7873[2], tmp7873[1], tmp7873[0]};
    assign tmp4549 = {tmp4548, const_408_0};
    assign tmp4561 = tmp3322 ^ tmp3554;
    assign tmp4566 = tmp4549 - tmp5532;
    assign tmp4567 = {tmp4566[8]};
    assign tmp4568 = {tmp4549[7]};
    assign tmp4569 = ~tmp4568;
    assign tmp4570 = tmp4567 ^ tmp4569;
    assign tmp4573 = tmp4570 ^ tmp171;
    assign tmp4574 = tmp4561 & tmp4573;
    assign tmp4583 = tmp5238 ^ tmp3554;
    assign tmp4591 = tmp5532 - tmp4549;
    assign tmp4592 = {tmp4591[8]};
    assign tmp4595 = tmp4592 ^ tmp171;
    assign tmp4598 = tmp4595 ^ tmp4569;
    assign tmp4599 = tmp5532 == tmp4549;
    assign tmp4600 = tmp4598 | tmp4599;
    assign tmp4601 = tmp3350 & tmp4600;
    assign tmp4602 = tmp4574 ? const_413_127 : tmp4549;
    assign tmp4603 = tmp4601 ? _ver_out_tmp_11 : tmp4602;
    assign tmp4606 = tmp7857 - tmp4603;
    assign tmp4607 = {tmp4606[8]};
    assign tmp4610 = tmp4607 ^ tmp3551;
    assign tmp4611 = {tmp4603[7]};
    assign tmp4612 = ~tmp4611;
    assign tmp4613 = tmp4610 ^ tmp4612;
    assign tmp4614 = tmp4547 & tmp4613;
    assign tmp4617 = tmp7877 - tmp7861;
    assign tmp4619 = {tmp7877[7]};
    assign tmp4621 = tmp3562 ^ tmp4246;
    assign tmp4623 = ~tmp5749;
    assign tmp4624 = tmp4621 ^ tmp4623;
    assign tmp4625 = tmp4614 & tmp4624;
    assign tmp4626 = {tmp7877[5], tmp7877[4], tmp7877[3], tmp7877[2], tmp7877[1], tmp7877[0]};
    assign tmp4627 = {tmp4626, const_415_0};
    assign tmp4633 = {tmp3970[8]};
    assign tmp4644 = tmp4627 - tmp5532;
    assign tmp4645 = {tmp4644[8]};
    assign tmp4646 = {tmp4627[7]};
    assign tmp4648 = tmp4645 ^ tmp4675;
    assign tmp4651 = tmp4648 ^ tmp171;
    assign tmp4652 = tmp5300 & tmp4651;
    assign tmp4669 = tmp5532 - tmp4627;
    assign tmp4670 = {tmp4669[8]};
    assign tmp4673 = tmp4670 ^ tmp171;
    assign tmp4675 = ~tmp4646;
    assign tmp4676 = tmp4673 ^ tmp4675;
    assign tmp4677 = tmp5532 == tmp4627;
    assign tmp4678 = tmp4676 | tmp4677;
    assign tmp4679 = tmp5325 & tmp4678;
    assign tmp4680 = tmp4652 ? const_420_127 : tmp4627;
    assign tmp4681 = tmp4679 ? _ver_out_tmp_12 : tmp4680;
    assign tmp4684 = tmp7861 - tmp4681;
    assign tmp4685 = {tmp4684[8]};
    assign tmp4688 = tmp4685 ^ tmp4623;
    assign tmp4689 = {tmp4681[7]};
    assign tmp4690 = ~tmp4689;
    assign tmp4691 = tmp4688 ^ tmp4690;
    assign tmp4692 = tmp4625 & tmp4691;
    assign tmp4698 = ~tmp3579;
    assign tmp4699 = tmp3575 ^ tmp4698;
    assign tmp4702 = tmp4699 ^ tmp4164;
    assign tmp4703 = tmp4692 & tmp4702;
    assign tmp4704 = {tmp7881[5], tmp7881[4], tmp7881[3], tmp7881[2], tmp7881[1], tmp7881[0]};
    assign tmp4705 = {tmp4704, const_422_0};
    assign tmp4711 = {tmp5374[8]};
    assign tmp4722 = tmp4705 - tmp5532;
    assign tmp4723 = {tmp4722[8]};
    assign tmp4724 = {tmp4705[7]};
    assign tmp4725 = ~tmp4724;
    assign tmp4726 = tmp4723 ^ tmp4725;
    assign tmp4729 = tmp4726 ^ tmp171;
    assign tmp4730 = tmp3473 & tmp4729;
    assign tmp4747 = tmp5532 - tmp4705;
    assign tmp4748 = {tmp4747[8]};
    assign tmp4751 = tmp4748 ^ tmp171;
    assign tmp4754 = tmp4751 ^ tmp4725;
    assign tmp4755 = tmp5532 == tmp4705;
    assign tmp4756 = tmp4754 | tmp4755;
    assign tmp4757 = tmp3498 & tmp4756;
    assign tmp4758 = tmp4730 ? const_427_127 : tmp4705;
    assign tmp4759 = tmp4757 ? _ver_out_tmp_15 : tmp4758;
    assign tmp4762 = tmp7865 - tmp4759;
    assign tmp4763 = {tmp4762[8]};
    assign tmp4766 = tmp4763 ^ tmp4164;
    assign tmp4767 = {tmp4759[7]};
    assign tmp4768 = ~tmp4767;
    assign tmp4769 = tmp4766 ^ tmp4768;
    assign tmp4770 = tmp4703 & tmp4769;
    assign tmp4817 = {tmp7853[7], tmp7853[6], tmp7853[5], tmp7853[4], tmp7853[3], tmp7853[2], tmp7853[1]};
    assign tmp4845 = {tmp7857[7], tmp7857[6], tmp7857[5], tmp7857[4], tmp7857[3], tmp7857[2], tmp7857[1]};
    assign tmp4874 = {tmp2948[6]};
    assign tmp4876 = {tmp4874, tmp2948};
    assign tmp4927 = tmp5045 & tmp4770;
    assign tmp4928 = tmp4927 & tmp7849;
    assign tmp4992 = ~tmp2981;
    assign tmp5018 = ~tmp3644;
    assign tmp5045 = tmp6670 & tmp5069;
    assign tmp5069 = ~tmp4259;
    assign tmp5074 = tmp4927 & tmp5447;
    assign tmp5136 = {tmp7869[7]};
    assign tmp5143 = tmp3239 - tmp5532;
    assign tmp5144 = {tmp5143[8]};
    assign tmp5146 = ~tmp3286;
    assign tmp5168 = tmp5532 - tmp3239;
    assign tmp5176 = tmp5532 == tmp3239;
    assign tmp5206 = {tmp7873[6], tmp7873[5], tmp7873[4], tmp7873[3], tmp7873[2], tmp7873[1], tmp7873[0]};
    assign tmp5207 = {tmp5206, const_438_0};
    assign tmp5226 = {tmp5207[7]};
    assign tmp5227 = ~tmp5226;
    assign tmp5228 = tmp5668 ^ tmp5227;
    assign tmp5229 = {tmp5532[7]};
    assign tmp5232 = tmp4561 & tmp5674;
    assign tmp5238 = {tmp5680[8]};
    assign tmp5259 = tmp3350 & tmp5701;
    assign tmp5287 = {tmp7877[6], tmp7877[5], tmp7877[4], tmp7877[3], tmp7877[2], tmp7877[1], tmp7877[0]};
    assign tmp5297 = tmp4633 ^ tmp171;
    assign tmp5300 = tmp5297 ^ tmp4246;
    assign tmp5306 = {tmp3404[8]};
    assign tmp5309 = tmp5306 ^ tmp3435;
    assign tmp5312 = tmp5309 ^ tmp171;
    assign tmp5313 = tmp5300 & tmp5312;
    assign tmp5325 = tmp3421 ^ tmp171;
    assign tmp5342 = tmp5836 ? _ver_out_tmp_25 : tmp3440;
    assign tmp5355 = tmp4311 & tmp7848;
    assign tmp5374 = tmp5532 - tmp7881;
    assign tmp5386 = tmp3461 - tmp5532;
    assign tmp5387 = {tmp5386[8]};
    assign tmp5388 = {tmp3461[7]};
    assign tmp5390 = tmp5387 ^ tmp5966;
    assign tmp5418 = tmp3507 ^ tmp5966;
    assign tmp5447 = ~tmp7849;
    assign tmp5449 = {tmp7853[6], tmp7853[5], tmp7853[4], tmp7853[3], tmp7853[2], tmp7853[1], tmp7853[0]};
    assign tmp5450 = {tmp5449, const_459_0};
    assign tmp5456 = {tmp6079[8]};
    assign tmp5462 = tmp6083 ^ tmp3762;
    assign tmp5467 = tmp5450 - tmp5532;
    assign tmp5468 = {tmp5467[8]};
    assign tmp5469 = {tmp5450[7]};
    assign tmp5470 = ~tmp5469;
    assign tmp5471 = tmp5468 ^ tmp5470;
    assign tmp5474 = tmp5471 ^ tmp171;
    assign tmp5475 = tmp5462 & tmp5474;
    assign tmp5484 = tmp3760 ^ tmp3762;
    assign tmp5487 = tmp5484 ^ tmp171;
    assign tmp5492 = tmp5532 - tmp5450;
    assign tmp5493 = {tmp5492[8]};
    assign tmp5496 = tmp5493 ^ tmp171;
    assign tmp5499 = tmp5496 ^ tmp5470;
    assign tmp5500 = tmp5532 == tmp5450;
    assign tmp5501 = tmp5499 | tmp5500;
    assign tmp5502 = tmp5487 & tmp5501;
    assign tmp5503 = tmp5475 ? const_464_127 : tmp5450;
    assign tmp5504 = tmp5502 ? _ver_out_tmp_30 : tmp5503;
    assign tmp5507 = tmp7869 - tmp5504;
    assign tmp5508 = {tmp5507[8]};
    assign tmp5510 = ~tmp5136;
    assign tmp5511 = tmp5508 ^ tmp5510;
    assign tmp5512 = {tmp5504[7]};
    assign tmp5513 = ~tmp5512;
    assign tmp5514 = tmp5511 ^ tmp5513;
    assign tmp5521 = tmp5532 - tmp7869;
    assign tmp5525 = tmp3245 ^ tmp171;
    assign tmp5528 = tmp5525 ^ tmp5510;
    assign tmp5532 = {tmp2736, const_468_0};
    assign tmp5540 = tmp3260 ^ tmp171;
    assign tmp5541 = tmp5528 & tmp5540;
    assign tmp5546 = tmp7869 - tmp5532;
    assign tmp5550 = tmp3270 ^ tmp5510;
    assign tmp5553 = tmp5550 ^ tmp171;
    assign tmp5569 = tmp5541 ? const_471_127 : tmp3239;
    assign tmp5570 = tmp3291 ? _ver_out_tmp_34 : tmp5569;
    assign tmp5573 = tmp7853 - tmp5570;
    assign tmp5574 = {tmp5573[8]};
    assign tmp5577 = tmp5574 ^ tmp3762;
    assign tmp5578 = {tmp5570[7]};
    assign tmp5579 = ~tmp5578;
    assign tmp5580 = tmp5577 ^ tmp5579;
    assign tmp5581 = tmp5514 & tmp5580;
    assign tmp5582 = {tmp7857[6], tmp7857[5], tmp7857[4], tmp7857[3], tmp7857[2], tmp7857[1], tmp7857[0]};
    assign tmp5583 = {tmp5582, const_473_0};
    assign tmp5595 = tmp3857 ^ tmp3551;
    assign tmp5600 = tmp5583 - tmp5532;
    assign tmp5601 = {tmp5600[8]};
    assign tmp5603 = ~tmp5630;
    assign tmp5604 = tmp5601 ^ tmp5603;
    assign tmp5607 = tmp5604 ^ tmp171;
    assign tmp5608 = tmp5595 & tmp5607;
    assign tmp5625 = tmp5532 - tmp5583;
    assign tmp5626 = {tmp5625[8]};
    assign tmp5629 = tmp5626 ^ tmp171;
    assign tmp5630 = {tmp5583[7]};
    assign tmp5632 = tmp5629 ^ tmp5603;
    assign tmp5633 = tmp5532 == tmp5583;
    assign tmp5634 = tmp5632 | tmp5633;
    assign tmp5635 = tmp6274 & tmp5634;
    assign tmp5636 = tmp5608 ? const_478_127 : tmp5583;
    assign tmp5637 = tmp5635 ? _ver_out_tmp_36 : tmp5636;
    assign tmp5640 = tmp7873 - tmp5637;
    assign tmp5641 = {tmp5640[8]};
    assign tmp5644 = tmp5641 ^ tmp3554;
    assign tmp5645 = {tmp5637[7]};
    assign tmp5646 = ~tmp5645;
    assign tmp5647 = tmp5644 ^ tmp5646;
    assign tmp5648 = tmp5581 & tmp5647;
    assign tmp5660 = {tmp7873[7]};
    assign tmp5667 = tmp5207 - tmp5532;
    assign tmp5668 = {tmp5667[8]};
    assign tmp5674 = tmp5228 ^ tmp171;
    assign tmp5680 = tmp7873 - tmp5532;
    assign tmp5692 = tmp5532 - tmp5207;
    assign tmp5693 = {tmp5692[8]};
    assign tmp5696 = tmp5693 ^ tmp171;
    assign tmp5699 = tmp5696 ^ tmp5227;
    assign tmp5700 = tmp5532 == tmp5207;
    assign tmp5701 = tmp5699 | tmp5700;
    assign tmp5707 = tmp7857 - tmp3367;
    assign tmp5708 = {tmp5707[8]};
    assign tmp5711 = tmp5708 ^ tmp3551;
    assign tmp5712 = {tmp3367[7]};
    assign tmp5713 = ~tmp5712;
    assign tmp5714 = tmp5711 ^ tmp5713;
    assign tmp5715 = tmp5648 & tmp5714;
    assign tmp5716 = {tmp7861[6], tmp7861[5], tmp7861[4], tmp7861[3], tmp7861[2], tmp7861[1], tmp7861[0]};
    assign tmp5717 = {tmp5716, const_487_0};
    assign tmp5722 = tmp5532 - tmp7861;
    assign tmp5723 = {tmp5722[8]};
    assign tmp5726 = tmp5723 ^ tmp171;
    assign tmp5734 = tmp5717 - tmp5532;
    assign tmp5735 = {tmp5734[8]};
    assign tmp5737 = ~tmp5764;
    assign tmp5738 = tmp5735 ^ tmp5737;
    assign tmp5741 = tmp5738 ^ tmp171;
    assign tmp5742 = tmp3994 & tmp5741;
    assign tmp5748 = {tmp6415[8]};
    assign tmp5749 = {tmp7861[7]};
    assign tmp5751 = tmp5748 ^ tmp4623;
    assign tmp5759 = tmp5532 - tmp5717;
    assign tmp5760 = {tmp5759[8]};
    assign tmp5763 = tmp5760 ^ tmp171;
    assign tmp5764 = {tmp5717[7]};
    assign tmp5766 = tmp5763 ^ tmp5737;
    assign tmp5767 = tmp5532 == tmp5717;
    assign tmp5768 = tmp5766 | tmp5767;
    assign tmp5769 = tmp6422 & tmp5768;
    assign tmp5770 = tmp5742 ? const_492_127 : tmp5717;
    assign tmp5771 = tmp5769 ? _ver_out_tmp_42 : tmp5770;
    assign tmp5774 = tmp7877 - tmp5771;
    assign tmp5775 = {tmp5774[8]};
    assign tmp5778 = tmp5775 ^ tmp4246;
    assign tmp5779 = {tmp5771[7]};
    assign tmp5780 = ~tmp5779;
    assign tmp5781 = tmp5778 ^ tmp5780;
    assign tmp5782 = tmp5715 & tmp5781;
    assign tmp5784 = {tmp5287, const_494_0};
    assign tmp5815 = {tmp3417[8]};
    assign tmp5831 = {tmp5784[7]};
    assign tmp5834 = tmp5532 == tmp5784;
    assign tmp5836 = tmp5325 & tmp3438;
    assign tmp5841 = tmp7861 - tmp5342;
    assign tmp5842 = {tmp5841[8]};
    assign tmp5845 = tmp5842 ^ tmp4623;
    assign tmp5846 = {tmp5342[7]};
    assign tmp5847 = ~tmp5846;
    assign tmp5848 = tmp5845 ^ tmp5847;
    assign tmp5849 = tmp5782 & tmp5848;
    assign tmp5850 = {tmp7865[6], tmp7865[5], tmp7865[4], tmp7865[3], tmp7865[2], tmp7865[1], tmp7865[0]};
    assign tmp5851 = {tmp5850, const_501_0};
    assign tmp5863 = tmp4125 ^ tmp4164;
    assign tmp5868 = tmp5851 - tmp5532;
    assign tmp5869 = {tmp5868[8]};
    assign tmp5871 = ~tmp5898;
    assign tmp5872 = tmp5869 ^ tmp5871;
    assign tmp5875 = tmp5872 ^ tmp171;
    assign tmp5876 = tmp5863 & tmp5875;
    assign tmp5881 = tmp7865 - tmp5532;
    assign tmp5882 = {tmp5881[8]};
    assign tmp5885 = tmp5882 ^ tmp4164;
    assign tmp5893 = tmp5532 - tmp5851;
    assign tmp5894 = {tmp5893[8]};
    assign tmp5897 = tmp5894 ^ tmp171;
    assign tmp5898 = {tmp5851[7]};
    assign tmp5900 = tmp5897 ^ tmp5871;
    assign tmp5901 = tmp5532 == tmp5851;
    assign tmp5902 = tmp5900 | tmp5901;
    assign tmp5903 = tmp6570 & tmp5902;
    assign tmp5904 = tmp5876 ? const_506_127 : tmp5851;
    assign tmp5905 = tmp5903 ? _ver_out_tmp_3 : tmp5904;
    assign tmp5908 = tmp7881 - tmp5905;
    assign tmp5909 = {tmp5908[8]};
    assign tmp5912 = tmp5909 ^ tmp4698;
    assign tmp5913 = {tmp5905[7]};
    assign tmp5914 = ~tmp5913;
    assign tmp5915 = tmp5912 ^ tmp5914;
    assign tmp5916 = tmp5849 & tmp5915;
    assign tmp5942 = tmp5390 ^ tmp171;
    assign tmp5960 = tmp5532 - tmp3461;
    assign tmp5966 = ~tmp5388;
    assign tmp5970 = tmp3498 & tmp3512;
    assign tmp5971 = tmp3486 ? const_513_127 : tmp3461;
    assign tmp5975 = tmp7865 - tmp3515;
    assign tmp5976 = {tmp5975[8]};
    assign tmp5979 = tmp5976 ^ tmp4164;
    assign tmp5980 = {tmp3515[7]};
    assign tmp5981 = ~tmp5980;
    assign tmp5982 = tmp5979 ^ tmp5981;
    assign tmp5983 = tmp5916 & tmp5982;
    assign tmp6058 = tmp6205 & tmp5983;
    assign tmp6067 = {tmp6084, tmp6084};
    assign tmp6074 = {tmp3713[7], tmp3713[6], tmp3713[5], tmp3713[4], tmp3713[3], tmp3713[2], tmp3713[1], tmp3713[0]};
    assign tmp6079 = tmp5532 - tmp7853;
    assign tmp6083 = tmp5456 ^ tmp171;
    assign tmp6084 = {tmp7853[7]};
    assign tmp6104 = tmp6074 - tmp5532;
    assign tmp6105 = {tmp6104[8]};
    assign tmp6111 = tmp3748 ^ tmp171;
    assign tmp6132 = {tmp3771[9]};
    assign tmp6138 = tmp3775 ^ tmp6538;
    assign tmp6139 = tmp5487 & tmp6138;
    assign tmp6144 = tmp5532 - tmp6074;
    assign tmp6145 = {tmp6144[8]};
    assign tmp6148 = tmp6145 ^ tmp171;
    assign tmp6151 = tmp6148 ^ tmp3747;
    assign tmp6153 = tmp6151 | tmp3752;
    assign tmp6156 = tmp3794 ? _ver_out_tmp_55 : tmp3795;
    assign tmp6205 = tmp5045 & tmp6623;
    assign tmp6210 = tmp5532 - tmp7873;
    assign tmp6211 = {const_534_0, const_534_0};
    assign tmp6213 = tmp3833 ? tmp2534 : tmp6210;
    assign tmp6221 = {tmp3846[9], tmp3846[8], tmp3846[7], tmp3846[6], tmp3846[5], tmp3846[4], tmp3846[3], tmp3846[2], tmp3846[1], tmp3846[0]};
    assign tmp6222 = {tmp6221[7], tmp6221[6], tmp6221[5], tmp6221[4], tmp6221[3], tmp6221[2], tmp6221[1], tmp6221[0]};
    assign tmp6240 = {tmp3865[9]};
    assign tmp6243 = tmp6240 ^ tmp6538;
    assign tmp6244 = {tmp6213[8]};
    assign tmp6245 = ~tmp6244;
    assign tmp6246 = tmp6243 ^ tmp6245;
    assign tmp6247 = tmp5595 & tmp6246;
    assign tmp6253 = {tmp3878[8]};
    assign tmp6256 = tmp6253 ^ tmp6298;
    assign tmp6259 = tmp6256 ^ tmp171;
    assign tmp6261 = tmp6259 | tmp6300;
    assign tmp6262 = tmp6247 & tmp6261;
    assign tmp6274 = tmp3897 ^ tmp171;
    assign tmp6279 = tmp6213 - tmp6533;
    assign tmp6283 = tmp3906 ^ tmp6245;
    assign tmp6286 = tmp6283 ^ tmp6538;
    assign tmp6287 = tmp6274 & tmp6286;
    assign tmp6292 = tmp5532 - tmp6222;
    assign tmp6293 = {tmp6292[8]};
    assign tmp6296 = tmp6293 ^ tmp171;
    assign tmp6297 = {tmp6222[7]};
    assign tmp6298 = ~tmp6297;
    assign tmp6300 = tmp5532 == tmp6222;
    assign tmp6303 = tmp6262 ? const_541_127 : tmp6222;
    assign tmp6304 = tmp3928 ? _ver_out_tmp_60 : tmp6303;
    assign tmp6355 = _ver_out_tmp_61 == tmp7877;
    assign tmp6368 = tmp3976 + tmp3979;
    assign tmp6369 = {tmp6368[9], tmp6368[8], tmp6368[7], tmp6368[6], tmp6368[5], tmp6368[4], tmp6368[3], tmp6368[2], tmp6368[1], tmp6368[0]};
    assign tmp6370 = {tmp6369[7], tmp6369[6], tmp6369[5], tmp6369[4], tmp6369[3], tmp6369[2], tmp6369[1], tmp6369[0]};
    assign tmp6384 = {const_549_0, const_549_0, const_549_0, const_549_0, const_549_0, const_549_0, const_549_0, const_549_0};
    assign tmp6388 = {tmp3999[9]};
    assign tmp6394 = tmp4003 ^ tmp4005;
    assign tmp6400 = tmp6370 - tmp5532;
    assign tmp6401 = {tmp6400[8]};
    assign tmp6402 = {tmp6370[7]};
    assign tmp6404 = tmp6401 ^ tmp6446;
    assign tmp6407 = tmp6404 ^ tmp171;
    assign tmp6410 = tmp4007 & tmp4021;
    assign tmp6415 = tmp7861 - tmp5532;
    assign tmp6422 = tmp5751 ^ tmp171;
    assign tmp6427 = tmp3973 - tmp6533;
    assign tmp6440 = tmp5532 - tmp6370;
    assign tmp6444 = tmp4053 ^ tmp171;
    assign tmp6446 = ~tmp6402;
    assign tmp6447 = tmp6444 ^ tmp6446;
    assign tmp6449 = tmp6447 | tmp4060;
    assign tmp6450 = tmp4047 & tmp6449;
    assign tmp6451 = tmp6410 ? const_554_127 : tmp6370;
    assign tmp6509 = tmp4101 ? tmp2534 : tmp5374;
    assign tmp6511 = {tmp4163, tmp4163};
    assign tmp6512 = {tmp6511, tmp7865};
    assign tmp6516 = tmp6512 + tmp4113;
    assign tmp6517 = {tmp6516[9], tmp6516[8], tmp6516[7], tmp6516[6], tmp6516[5], tmp6516[4], tmp6516[3], tmp6516[2], tmp6516[1], tmp6516[0]};
    assign tmp6533 = {tmp6384, const_562_0};
    assign tmp6535 = tmp6533 - tmp6509;
    assign tmp6537 = {tmp6533[8]};
    assign tmp6538 = ~tmp6537;
    assign tmp6539 = tmp4134 ^ tmp6538;
    assign tmp6541 = ~tmp6577;
    assign tmp6542 = tmp6539 ^ tmp6541;
    assign tmp6543 = tmp5863 & tmp6542;
    assign tmp6552 = tmp4147 ^ tmp4149;
    assign tmp6555 = tmp6552 ^ tmp171;
    assign tmp6557 = tmp6555 | tmp4194;
    assign tmp6558 = tmp6543 & tmp6557;
    assign tmp6570 = tmp5885 ^ tmp171;
    assign tmp6575 = tmp6509 - tmp6533;
    assign tmp6577 = {tmp6509[8]};
    assign tmp6579 = tmp4174 ^ tmp6541;
    assign tmp6583 = tmp6570 & tmp4180;
    assign tmp6588 = tmp5532 - tmp4116;
    assign tmp6592 = tmp4187 ^ tmp171;
    assign tmp6595 = tmp6592 ^ tmp4149;
    assign tmp6597 = tmp6595 | tmp4194;
    assign tmp6598 = tmp6583 & tmp6597;
    assign tmp6599 = tmp6558 ? const_567_127 : tmp4116;
    assign tmp6623 = ~tmp4770;
    assign tmp6651 = tmp6205 & tmp6676;
    assign tmp6670 = tmp4456 & tmp5018;
    assign tmp6676 = ~tmp5983;
    assign tmp6725 = tmp520 == const_573_1;
    assign tmp6734 = {const_579_0, tmp11};
    assign tmp6735 = tmp6725 ? tmp2459 : tmp6734;
    assign tmp6744 = tmp7041 ? tmp2534 : tmp7321;
    assign tmp6746 = {const_586_0, tmp15};
    assign tmp6747 = tmp7040 ? tmp6744 : tmp6746;
    assign tmp6750 = tmp6735 - tmp6747;
    assign tmp6751 = {tmp6750[9]};
    assign tmp6752 = {tmp6735[8]};
    assign tmp6753 = ~tmp6752;
    assign tmp6754 = tmp6751 ^ tmp6753;
    assign tmp6755 = {tmp6747[8]};
    assign tmp6756 = ~tmp6755;
    assign tmp6757 = tmp6754 ^ tmp6756;
    assign tmp6759 = tmp1615 == const_587_1;
    assign tmp6763 = tmp5532 - tmp12;
    assign tmp6766 = tmp1030 ? tmp2534 : tmp6763;
    assign tmp6769 = tmp6759 ? tmp6766 : tmp7074;
    assign tmp6771 = tmp938 == const_594_1;
    assign tmp6780 = {const_600_0, tmp16};
    assign tmp6781 = tmp6771 ? tmp7088 : tmp6780;
    assign tmp6784 = tmp6769 - tmp6781;
    assign tmp6785 = {tmp6784[9]};
    assign tmp6786 = {tmp6769[8]};
    assign tmp6787 = ~tmp6786;
    assign tmp6788 = tmp6785 ^ tmp6787;
    assign tmp6789 = {tmp6781[8]};
    assign tmp6790 = ~tmp6789;
    assign tmp6791 = tmp6788 ^ tmp6790;
    assign tmp6792 = tmp6757 & tmp6791;
    assign tmp6803 = {const_607_0, tmp13};
    assign tmp6807 = tmp17 == _ver_out_tmp_82;
    assign tmp6813 = tmp6807 ? tmp2534 : tmp1973;
    assign tmp6819 = tmp7116 - tmp7132;
    assign tmp6820 = {tmp6819[9]};
    assign tmp6821 = {tmp7116[8]};
    assign tmp6822 = ~tmp6821;
    assign tmp6823 = tmp6820 ^ tmp6822;
    assign tmp6825 = ~tmp7140;
    assign tmp6826 = tmp6823 ^ tmp6825;
    assign tmp6827 = tmp6792 & tmp6826;
    assign tmp6829 = tmp644 == const_615_1;
    assign tmp6830 = tmp14 == _ver_out_tmp_84;
    assign tmp6838 = {const_621_0, tmp14};
    assign tmp6839 = tmp6829 ? tmp2516 : tmp6838;
    assign tmp6841 = tmp7162 == const_622_1;
    assign tmp6845 = tmp5532 - tmp18;
    assign tmp6848 = tmp2586 ? tmp2534 : tmp6845;
    assign tmp6854 = tmp6839 - tmp7173;
    assign tmp6855 = {tmp6854[9]};
    assign tmp6856 = {tmp6839[8]};
    assign tmp6857 = ~tmp6856;
    assign tmp6858 = tmp6855 ^ tmp6857;
    assign tmp6859 = {tmp7173[8]};
    assign tmp6861 = tmp6858 ^ tmp7182;
    assign tmp6862 = tmp6827 & tmp6861;
    assign tmp6958 = tmp6972 & tmp6862;
    assign tmp6972 = tmp4311 & tmp7383;
    assign tmp7035 = {tmp6735[8], tmp6735[7], tmp6735[6], tmp6735[5], tmp6735[4], tmp6735[3], tmp6735[2], tmp6735[1]};
    assign tmp7036 = {tmp7035[7]};
    assign tmp7038 = {tmp7036, tmp7035};
    assign tmp7040 = tmp2623 == const_638_1;
    assign tmp7041 = tmp15 == _ver_out_tmp_33;
    assign tmp7053 = tmp6747 - tmp7038;
    assign tmp7054 = {tmp7053[9]};
    assign tmp7055 = {tmp7038[8]};
    assign tmp7056 = ~tmp7055;
    assign tmp7057 = tmp7054 ^ tmp7056;
    assign tmp7060 = tmp7057 ^ tmp6756;
    assign tmp7061 = tmp7038 == tmp6747;
    assign tmp7062 = tmp7060 | tmp7061;
    assign tmp7063 = tmp19 & tmp7062;
    assign tmp7074 = {const_651_0, tmp12};
    assign tmp7076 = {tmp6769[8], tmp6769[7], tmp6769[6], tmp6769[5], tmp6769[4], tmp6769[3], tmp6769[2], tmp6769[1]};
    assign tmp7077 = {tmp7076[7]};
    assign tmp7079 = {tmp7077, tmp7076};
    assign tmp7088 = tmp2548 ? tmp2534 : tmp1860;
    assign tmp7094 = tmp6781 - tmp7079;
    assign tmp7095 = {tmp7094[9]};
    assign tmp7096 = {tmp7079[8]};
    assign tmp7097 = ~tmp7096;
    assign tmp7098 = tmp7095 ^ tmp7097;
    assign tmp7101 = tmp7098 ^ tmp6790;
    assign tmp7102 = tmp7079 == tmp6781;
    assign tmp7103 = tmp7101 | tmp7102;
    assign tmp7104 = tmp7063 & tmp7103;
    assign tmp7106 = tmp550 == const_659_1;
    assign tmp7116 = tmp7106 ? tmp2877 : tmp6803;
    assign tmp7117 = {tmp7116[8], tmp7116[7], tmp7116[6], tmp7116[5], tmp7116[4], tmp7116[3], tmp7116[2], tmp7116[1]};
    assign tmp7118 = {tmp7117[7]};
    assign tmp7120 = {tmp7118, tmp7117};
    assign tmp7121 = {tmp17[7]};
    assign tmp7122 = tmp7121 == const_666_1;
    assign tmp7131 = {const_672_0, tmp17};
    assign tmp7132 = tmp7122 ? tmp6813 : tmp7131;
    assign tmp7135 = tmp7132 - tmp7120;
    assign tmp7136 = {tmp7135[9]};
    assign tmp7137 = {tmp7120[8]};
    assign tmp7138 = ~tmp7137;
    assign tmp7139 = tmp7136 ^ tmp7138;
    assign tmp7140 = {tmp7132[8]};
    assign tmp7142 = tmp7139 ^ tmp6825;
    assign tmp7143 = tmp7120 == tmp7132;
    assign tmp7144 = tmp7142 | tmp7143;
    assign tmp7145 = tmp7104 & tmp7144;
    assign tmp7158 = {tmp6839[8], tmp6839[7], tmp6839[6], tmp6839[5], tmp6839[4], tmp6839[3], tmp6839[2], tmp6839[1]};
    assign tmp7159 = {tmp7158[7]};
    assign tmp7161 = {tmp7159, tmp7158};
    assign tmp7162 = {tmp18[7]};
    assign tmp7172 = {const_686_0, tmp18};
    assign tmp7173 = tmp6841 ? tmp6848 : tmp7172;
    assign tmp7176 = tmp7173 - tmp7161;
    assign tmp7177 = {tmp7176[9]};
    assign tmp7178 = {tmp7161[8]};
    assign tmp7179 = ~tmp7178;
    assign tmp7180 = tmp7177 ^ tmp7179;
    assign tmp7182 = ~tmp6859;
    assign tmp7183 = tmp7180 ^ tmp7182;
    assign tmp7184 = tmp7161 == tmp7173;
    assign tmp7185 = tmp7183 | tmp7184;
    assign tmp7186 = tmp7145 & tmp7185;
    assign tmp7223 = {tmp11[7], tmp11[6], tmp11[5], tmp11[4], tmp11[3], tmp11[2], tmp11[1]};
    assign tmp7224 = {tmp7223[6]};
    assign tmp7226 = {tmp7224, tmp7223};
    assign tmp7242 = ~tmp6862;
    assign tmp7243 = tmp6972 & tmp7242;
    assign tmp7244 = tmp7243 & tmp7186;
    assign tmp7246 = {tmp12[7], tmp12[6], tmp12[5], tmp12[4], tmp12[3], tmp12[2], tmp12[1]};
    assign tmp7247 = {tmp7246[6]};
    assign tmp7249 = {tmp7247, tmp7246};
    assign tmp7268 = tmp7244 & tmp7849;
    assign tmp7269 = {tmp13[7], tmp13[6], tmp13[5], tmp13[4], tmp13[3], tmp13[2], tmp13[1]};
    assign tmp7270 = {tmp7269[6]};
    assign tmp7272 = {tmp7270, tmp7269};
    assign tmp7292 = {tmp14[7], tmp14[6], tmp14[5], tmp14[4], tmp14[3], tmp14[2], tmp14[1]};
    assign tmp7293 = {tmp7292[6]};
    assign tmp7295 = {tmp7293, tmp7292};
    assign tmp7316 = {tmp268, const_689_0};
    assign tmp7321 = tmp5532 - tmp15;
    assign tmp7325 = tmp1320 ^ tmp171;
    assign tmp7327 = ~tmp2623;
    assign tmp7341 = tmp1326 & tmp1338;
    assign tmp7358 = tmp5532 - tmp7316;
    assign tmp7362 = tmp312 ^ tmp171;
    assign tmp7366 = tmp5532 == tmp7316;
    assign tmp7368 = tmp2628 & tmp320;
    assign tmp7370 = tmp7368 ? _ver_out_tmp_66 : tmp1367;
    assign tmp7383 = ~tmp7848;
    assign tmp7391 = {tmp16[6], tmp16[5], tmp16[4], tmp16[3], tmp16[2], tmp16[1], tmp16[0]};
    assign tmp7392 = {tmp7391, const_696_0};
    assign tmp7404 = tmp345 ^ tmp902;
    assign tmp7409 = tmp7392 - tmp5532;
    assign tmp7411 = {tmp7392[7]};
    assign tmp7412 = ~tmp7411;
    assign tmp7413 = tmp354 ^ tmp7412;
    assign tmp7416 = tmp7413 ^ tmp171;
    assign tmp7417 = tmp7404 & tmp7416;
    assign tmp7422 = tmp16 - tmp5532;
    assign tmp7434 = tmp5532 - tmp7392;
    assign tmp7435 = {tmp7434[8]};
    assign tmp7438 = tmp7435 ^ tmp171;
    assign tmp7441 = tmp7438 ^ tmp7412;
    assign tmp7442 = tmp5532 == tmp7392;
    assign tmp7443 = tmp7441 | tmp7442;
    assign tmp7445 = tmp7417 ? const_701_127 : tmp7392;
    assign tmp7446 = tmp388 ? _ver_out_tmp_68 : tmp7445;
    assign tmp7466 = tmp7244 & tmp5447;
    assign tmp7467 = {tmp17[6], tmp17[5], tmp17[4], tmp17[3], tmp17[2], tmp17[1], tmp17[0]};
    assign tmp7468 = {tmp7467, const_703_0};
    assign tmp7474 = {tmp1973[8]};
    assign tmp7486 = {tmp1400[8]};
    assign tmp7487 = {tmp7468[7]};
    assign tmp7488 = ~tmp7487;
    assign tmp7493 = tmp1980 & tmp1407;
    assign tmp7502 = tmp2014 ^ tmp1979;
    assign tmp7517 = tmp1429 ^ tmp7488;
    assign tmp7518 = tmp5532 == tmp7468;
    assign tmp7543 = {tmp18[6], tmp18[5], tmp18[4], tmp18[3], tmp18[2], tmp18[1], tmp18[0]};
    assign tmp7544 = {tmp7543, const_710_0};
    assign tmp7556 = tmp912 ^ tmp2354;
    assign tmp7561 = tmp7544 - tmp5532;
    assign tmp7562 = {tmp7561[8]};
    assign tmp7563 = {tmp7544[7]};
    assign tmp7565 = tmp7562 ^ tmp7592;
    assign tmp7568 = tmp7565 ^ tmp171;
    assign tmp7569 = tmp7556 & tmp7568;
    assign tmp7586 = tmp5532 - tmp7544;
    assign tmp7587 = {tmp7586[8]};
    assign tmp7590 = tmp7587 ^ tmp171;
    assign tmp7592 = ~tmp7563;
    assign tmp7593 = tmp7590 ^ tmp7592;
    assign tmp7594 = tmp5532 == tmp7544;
    assign tmp7595 = tmp7593 | tmp7594;
    assign tmp7596 = tmp2032 & tmp7595;
    assign tmp7597 = tmp7569 ? const_715_127 : tmp7544;
    assign tmp7598 = tmp7596 ? _ver_out_tmp_70 : tmp7597;
    assign tmp7636 = ~tmp7186;
    assign tmp7637 = tmp7243 & tmp7636;
    assign tmp7644 = tmp3298 & tmp2702;
    assign tmp7689 = tmp61 ? const_6_0 : tmp11;
    assign tmp7690 = tmp334 ? tmp1230 : tmp7689;
    assign tmp7691 = tmp421 ? tmp13 : tmp7690;
    assign tmp7692 = tmp988 ? tmp610 : tmp7691;
    assign tmp7693 = tmp1104 ? tmp2460 : tmp7692;
    assign tmp7694 = tmp1381 ? tmp1230 : tmp7693;
    assign tmp7695 = tmp1577 ? tmp12 : tmp7694;
    assign tmp7696 = tmp1709 ? tmp1675 : tmp7695;
    assign tmp7697 = tmp2193 ? tmp2460 : tmp7696;
    assign tmp7698 = tmp2892 ? tmp2460 : tmp7697;
    assign tmp7699 = tmp3055 ? tmp3588 : tmp7698;
    assign tmp7700 = tmp3201 ? tmp7853 : tmp7699;
    assign tmp7701 = tmp3698 ? tmp7869 : tmp7700;
    assign tmp7702 = tmp4359 ? tmp7869 : tmp7701;
    assign tmp7703 = tmp4928 ? tmp3588 : tmp7702;
    assign tmp7704 = tmp5074 ? tmp7853 : tmp7703;
    assign tmp7705 = tmp6058 ? tmp7869 : tmp7704;
    assign tmp7706 = tmp6958 ? tmp15 : tmp7705;
    assign tmp7707 = tmp7268 ? tmp7226 : tmp7706;
    assign tmp7708 = tmp61 ? const_7_2 : tmp12;
    assign tmp7709 = tmp334 ? tmp256 : tmp7708;
    assign tmp7710 = tmp421 ? tmp14 : tmp7709;
    assign tmp7711 = tmp988 ? tmp731 : tmp7710;
    assign tmp7712 = tmp1104 ? tmp2856 : tmp7711;
    assign tmp7713 = tmp1141 ? tmp11 : tmp7712;
    assign tmp7714 = tmp1577 ? tmp11 : tmp7713;
    assign tmp7715 = tmp1709 ? tmp11 : tmp7714;
    assign tmp7716 = tmp2892 ? tmp2856 : tmp7715;
    assign tmp7717 = tmp3055 ? tmp3038 : tmp7716;
    assign tmp7718 = tmp3201 ? tmp7857 : tmp7717;
    assign tmp7719 = tmp3698 ? tmp7873 : tmp7718;
    assign tmp7720 = tmp4359 ? tmp7873 : tmp7719;
    assign tmp7721 = tmp4928 ? tmp3038 : tmp7720;
    assign tmp7722 = tmp5074 ? tmp7857 : tmp7721;
    assign tmp7723 = tmp6058 ? tmp7873 : tmp7722;
    assign tmp7724 = tmp6958 ? tmp16 : tmp7723;
    assign tmp7725 = tmp7268 ? tmp7249 : tmp7724;
    assign tmp7726 = tmp61 ? const_8_1 : tmp13;
    assign tmp7727 = tmp122 ? tmp11 : tmp7726;
    assign tmp7728 = tmp421 ? tmp11 : tmp7727;
    assign tmp7729 = tmp988 ? tmp11 : tmp7728;
    assign tmp7730 = tmp1381 ? tmp1299 : tmp7729;
    assign tmp7731 = tmp1577 ? tmp14 : tmp7730;
    assign tmp7732 = tmp1709 ? tmp1800 : tmp7731;
    assign tmp7733 = tmp2193 ? tmp2120 : tmp7732;
    assign tmp7734 = tmp2892 ? tmp2120 : tmp7733;
    assign tmp7735 = tmp3055 ? tmp4876 : tmp7734;
    assign tmp7736 = tmp3201 ? tmp7861 : tmp7735;
    assign tmp7737 = tmp3698 ? tmp7877 : tmp7736;
    assign tmp7738 = tmp4359 ? tmp7877 : tmp7737;
    assign tmp7739 = tmp4928 ? tmp4876 : tmp7738;
    assign tmp7740 = tmp5074 ? tmp7861 : tmp7739;
    assign tmp7741 = tmp6058 ? tmp7877 : tmp7740;
    assign tmp7742 = tmp6958 ? tmp17 : tmp7741;
    assign tmp7743 = tmp7268 ? tmp7272 : tmp7742;
    assign tmp7744 = tmp61 ? const_9_0 : tmp14;
    assign tmp7745 = tmp122 ? tmp12 : tmp7744;
    assign tmp7746 = tmp421 ? tmp12 : tmp7745;
    assign tmp7747 = tmp988 ? tmp12 : tmp7746;
    assign tmp7748 = tmp1141 ? tmp13 : tmp7747;
    assign tmp7749 = tmp1577 ? tmp13 : tmp7748;
    assign tmp7750 = tmp1709 ? tmp13 : tmp7749;
    assign tmp7751 = tmp2892 ? tmp2517 : tmp7750;
    assign tmp7752 = tmp3055 ? tmp3633 : tmp7751;
    assign tmp7753 = tmp3201 ? tmp7865 : tmp7752;
    assign tmp7754 = tmp3698 ? tmp7881 : tmp7753;
    assign tmp7755 = tmp4359 ? tmp7881 : tmp7754;
    assign tmp7756 = tmp4928 ? tmp3633 : tmp7755;
    assign tmp7757 = tmp5074 ? tmp7865 : tmp7756;
    assign tmp7758 = tmp6058 ? tmp7881 : tmp7757;
    assign tmp7759 = tmp6958 ? tmp18 : tmp7758;
    assign tmp7760 = tmp7268 ? tmp7295 : tmp7759;
    assign tmp7761 = tmp61 ? const_10_0 : tmp15;
    assign tmp7762 = tmp334 ? tmp7370 : tmp7761;
    assign tmp7763 = tmp421 ? tmp17 : tmp7762;
    assign tmp7764 = tmp988 ? tmp852 : tmp7763;
    assign tmp7765 = tmp1104 ? tmp1062 : tmp7764;
    assign tmp7766 = tmp1381 ? tmp7370 : tmp7765;
    assign tmp7767 = tmp1577 ? tmp16 : tmp7766;
    assign tmp7768 = tmp1709 ? tmp1925 : tmp7767;
    assign tmp7769 = tmp2193 ? tmp1062 : tmp7768;
    assign tmp7770 = tmp3055 ? tmp7869 : tmp7769;
    assign tmp7771 = tmp3201 ? tmp5570 : tmp7770;
    assign tmp7772 = tmp3698 ? tmp6156 : tmp7771;
    assign tmp7773 = tmp4359 ? tmp7853 : tmp7772;
    assign tmp7774 = tmp4928 ? tmp7869 : tmp7773;
    assign tmp7775 = tmp5074 ? tmp5570 : tmp7774;
    assign tmp7776 = tmp6058 ? tmp6156 : tmp7775;
    assign tmp7777 = tmp6958 ? tmp11 : tmp7776;
    assign tmp7778 = tmp7466 ? tmp7370 : tmp7777;
    assign tmp7779 = tmp61 ? const_11_0 : tmp16;
    assign tmp7780 = tmp334 ? tmp7446 : tmp7779;
    assign tmp7781 = tmp421 ? tmp18 : tmp7780;
    assign tmp7782 = tmp988 ? tmp973 : tmp7781;
    assign tmp7783 = tmp1104 ? tmp2555 : tmp7782;
    assign tmp7784 = tmp1141 ? tmp15 : tmp7783;
    assign tmp7785 = tmp1577 ? tmp15 : tmp7784;
    assign tmp7786 = tmp1709 ? tmp15 : tmp7785;
    assign tmp7787 = tmp3055 ? tmp7873 : tmp7786;
    assign tmp7788 = tmp3201 ? tmp3367 : tmp7787;
    assign tmp7789 = tmp3698 ? tmp6304 : tmp7788;
    assign tmp7790 = tmp4359 ? tmp7857 : tmp7789;
    assign tmp7791 = tmp4928 ? tmp7873 : tmp7790;
    assign tmp7792 = tmp5074 ? tmp3367 : tmp7791;
    assign tmp7793 = tmp6058 ? tmp6304 : tmp7792;
    assign tmp7794 = tmp6958 ? tmp12 : tmp7793;
    assign tmp7795 = tmp7466 ? tmp7446 : tmp7794;
    assign tmp7796 = tmp61 ? const_12_0 : tmp17;
    assign tmp7797 = tmp122 ? tmp15 : tmp7796;
    assign tmp7798 = tmp421 ? tmp15 : tmp7797;
    assign tmp7799 = tmp988 ? tmp15 : tmp7798;
    assign tmp7800 = tmp1381 ? tmp1437 : tmp7799;
    assign tmp7801 = tmp1577 ? tmp18 : tmp7800;
    assign tmp7802 = tmp1709 ? tmp2050 : tmp7801;
    assign tmp7803 = tmp2193 ? tmp2174 : tmp7802;
    assign tmp7804 = tmp3055 ? tmp7877 : tmp7803;
    assign tmp7805 = tmp3201 ? tmp5342 : tmp7804;
    assign tmp7806 = tmp3698 ? tmp4064 : tmp7805;
    assign tmp7807 = tmp4359 ? tmp7861 : tmp7806;
    assign tmp7808 = tmp4928 ? tmp7877 : tmp7807;
    assign tmp7809 = tmp5074 ? tmp5342 : tmp7808;
    assign tmp7810 = tmp6058 ? tmp4064 : tmp7809;
    assign tmp7811 = tmp6958 ? tmp13 : tmp7810;
    assign tmp7812 = tmp7466 ? tmp1437 : tmp7811;
    assign tmp7813 = tmp61 ? const_13_1 : tmp18;
    assign tmp7814 = tmp122 ? tmp16 : tmp7813;
    assign tmp7815 = tmp421 ? tmp16 : tmp7814;
    assign tmp7816 = tmp988 ? tmp16 : tmp7815;
    assign tmp7817 = tmp1141 ? tmp17 : tmp7816;
    assign tmp7818 = tmp1577 ? tmp17 : tmp7817;
    assign tmp7819 = tmp1709 ? tmp17 : tmp7818;
    assign tmp7820 = tmp3055 ? tmp7881 : tmp7819;
    assign tmp7821 = tmp3201 ? tmp3515 : tmp7820;
    assign tmp7822 = tmp3698 ? tmp4198 : tmp7821;
    assign tmp7823 = tmp4359 ? tmp7865 : tmp7822;
    assign tmp7824 = tmp4928 ? tmp7881 : tmp7823;
    assign tmp7825 = tmp5074 ? tmp3515 : tmp7824;
    assign tmp7826 = tmp6058 ? tmp4198 : tmp7825;
    assign tmp7827 = tmp6958 ? tmp14 : tmp7826;
    assign tmp7828 = tmp7466 ? tmp7598 : tmp7827;
    assign tmp7829 = tmp61 ? const_14_0 : tmp19;
    assign tmp7830 = tmp1093 ? tmp19 : tmp7829;
    assign tmp7831 = tmp1127 ? tmp19 : tmp7830;
    assign tmp7832 = tmp2772 ? const_290_0 : tmp7831;
    assign tmp7833 = tmp2892 ? const_294_0 : tmp7832;
    assign tmp7834 = tmp3113 ? const_316_0 : tmp7833;
    assign tmp7835 = tmp3698 ? const_346_0 : tmp7834;
    assign tmp7836 = tmp4359 ? const_400_0 : tmp7835;
    assign tmp7837 = tmp4927 ? const_430_0 : tmp7836;
    assign tmp7838 = tmp6058 ? const_516_1 : tmp7837;
    assign tmp7839 = tmp6651 ? const_570_0 : tmp7838;
    assign tmp7840 = const_781_0 ? const_572_0 : tmp7839;
    assign tmp7841 = tmp6958 ? const_630_1 : tmp7840;
    assign tmp7842 = tmp7244 ? const_688_1 : tmp7841;
    assign tmp7843 = tmp7637 ? tmp19 : tmp7842;
    assign tmp7844 = const_780_0 ? tmp19 : tmp7843;
    assign tmp7845 = tmp2706 ? tmp2273 : const_719_0;
    assign tmp7846 = tmp2706 ? tmp2360 : const_720_0;
    assign tmp7847 = tmp2706 ? tmp2385 : const_721_0;
    assign tmp7848 = tmp2706 ? tmp2398 : const_722_0;
    assign tmp7849 = tmp2706 ? tmp2416 : const_723_0;
    assign tmp7852 = tmp2566 ? tmp2460 : tmp5532;
    assign tmp7853 = tmp2735 ? tmp11 : tmp7852;
    assign tmp7856 = tmp2566 ? tmp2856 : tmp5532;
    assign tmp7857 = tmp2735 ? tmp12 : tmp7856;
    assign tmp7860 = tmp2566 ? tmp2120 : tmp5532;
    assign tmp7861 = tmp2735 ? tmp13 : tmp7860;
    assign tmp7864 = tmp2566 ? tmp2517 : tmp5532;
    assign tmp7865 = tmp2735 ? tmp14 : tmp7864;
    assign tmp7868 = tmp2566 ? tmp1062 : tmp5532;
    assign tmp7869 = tmp2735 ? tmp15 : tmp7868;
    assign tmp7872 = tmp2566 ? tmp2555 : tmp5532;
    assign tmp7873 = tmp2735 ? tmp16 : tmp7872;
    assign tmp7876 = tmp2566 ? tmp2174 : tmp5532;
    assign tmp7877 = tmp2735 ? tmp17 : tmp7876;
    assign tmp7880 = tmp2566 ? tmp2593 : tmp5532;
    assign tmp7881 = tmp2735 ? tmp18 : tmp7880;
    assign tmp7882 = tmp2772 ? const_289_15 : my_calculator_out_z;
    assign tmp7883 = tmp2892 ? const_293_8 : tmp7882;
    assign tmp7884 = tmp3113 ? const_315_1 : tmp7883;
    assign tmp7885 = tmp3698 ? const_345_4 : tmp7884;
    assign tmp7886 = tmp4359 ? const_399_6 : tmp7885;
    assign tmp7887 = tmp4927 ? const_429_2 : tmp7886;
    assign tmp7888 = tmp6058 ? const_515_5 : tmp7887;
    assign tmp7889 = tmp6651 ? const_569_0 : tmp7888;
    assign tmp7890 = const_779_0 ? const_571_0 : tmp7889;
    assign tmp7891 = tmp6958 ? const_629_7 : tmp7890;
    assign tmp7892 = tmp7244 ? const_687_3 : tmp7891;
    assign tmp7893 = tmp7637 ? const_717_0 : tmp7892;
    assign tmp7894 = const_778_0 ? const_718_0 : tmp7893;
    assign tmp7902 = tmp7899 == tmp1165;
    assign tmp7904 = {tmp6211, const_742_2};
    assign tmp7905 = tmp7899 == tmp7904;
    assign tmp7906 = tmp7902 | tmp7905;
    assign tmp7908 = {tmp6211, const_744_3};
    assign tmp7909 = tmp7899 == tmp7908;
    assign tmp7910 = tmp7906 | tmp7909;
    assign tmp7912 = tmp7910 | tmp7939;
    assign tmp7915 = tmp7899 == tmp514;
    assign tmp7917 = {const_750_0, const_749_5};
    assign tmp7918 = tmp7899 == tmp7917;
    assign tmp7919 = tmp7915 | tmp7918;
    assign tmp7923 = tmp7919 | tmp7933;
    assign tmp7926 = tmp7899 == tmp1455;
    assign tmp7927 = tmp7923 | tmp7926;
    assign tmp7929 = tmp7927 | tmp7939;
    assign tmp7930 = tmp7899 == const_756_8;
    assign tmp7933 = tmp7899 == tmp1452;
    assign tmp7934 = tmp7930 | tmp7933;
    assign tmp7938 = tmp7934 | tmp7926;
    assign tmp7939 = tmp7899 == const_761_15;
    assign tmp7940 = tmp7938 | tmp7939;
    assign tmp7944 = {const_763_0, const_763_0, const_763_0, const_763_0};
    assign tmp7945 = {tmp7944, const_762_1};
    assign tmp7946 = tmp7895 + tmp7945;
    assign tmp7947 = {tmp7946[4], tmp7946[3], tmp7946[2], tmp7946[1], tmp7946[0]};
    assign tmp7949 = tmp7941 == const_764_4;
    assign tmp7950 = tmp7 & tmp7949;
    assign tmp7953 = tmp7941 == tmp75;
    assign tmp7954 = ~tmp7949;
    assign tmp7956 = tmp7961 & tmp7953;
    assign tmp7959 = tmp7941 == tmp1106;
    assign tmp7961 = tmp7 & tmp7954;
    assign tmp7962 = ~tmp7953;
    assign tmp7963 = tmp7961 & tmp7962;
    assign tmp7964 = tmp7963 & tmp7959;
    assign tmp7967 = tmp7941 == tmp2195;
    assign tmp7972 = ~tmp7959;
    assign tmp7973 = tmp7963 & tmp7972;
    assign tmp7974 = tmp7973 & tmp7967;
    assign tmp7975 = tmp7 ? tmp7947 : tmp7895;
    assign tmp7976 = tmp7950 ? const_765_8 : tmp7899;
    assign tmp7977 = tmp7956 ? my_calculator_out_z : tmp7976;
    assign tmp7978 = tmp7964 ? const_770_6 : tmp7977;
    assign tmp7979 = tmp7974 ? const_773_6 : tmp7978;

    // Registers
    always @(posedge clk)
    begin
        begin
            my_calculator_ctrl <= tmp7941;
            my_calculator_in_x <= tmp7942;
            my_calculator_in_y <= tmp7943;
            my_calculator_out_z <= tmp7894;
            tmp0 <= tmp4;
            tmp5 <= tmp8;
            tmp7 <= tmp10;
            tmp11 <= tmp7707;
            tmp12 <= tmp7725;
            tmp13 <= tmp7743;
            tmp14 <= tmp7760;
            tmp15 <= tmp7778;
            tmp16 <= tmp7795;
            tmp17 <= tmp7812;
            tmp18 <= tmp7828;
            tmp19 <= tmp7844;
            tmp7895 <= tmp7975;
            tmp7899 <= tmp7979;
        end
    end

    // Memory mem_0: tmp7896
    assign tmp7941 = mem_0[tmp7895];

    // Memory mem_1: tmp7897
    assign tmp7942 = mem_1[tmp7895];

    // Memory mem_2: tmp7898
    assign tmp7943 = mem_2[tmp7895];

endmodule

