// Simple tri-colour LED blink example.

// Correctly map pins for the iCE40UP5K SB_RGBA_DRV hard macro.

`define GREENPWM RGB0PWM
`define REDPWM   RGB1PWM
`define BLUEPWM  RGB2PWM

// taken (mostly) from
// https://github.com/im-tomu/fomu-workshop/blob/master/hdl/verilog/blink-expanded/blink.v

module top (
    // 48MHz Clock input
    // --------
    input clki,
    // LED outputs
    // --------
    output rgb0,
    output rgb1,
    output rgb2,
    // User touchable pins
    // --------
    // Connect 1-2 to enable blue LED
    input  user_1,
    output user_2,
    // Connect 3-4 to enable red LED
    output user_3,
    input  user_4,
    // USB Pins (which should be statically driven if not being used).
    // --------
    output usb_dp,
    output usb_dn,
    output usb_dp_pu
);

    // Assign USB pins to "0" so as to disconnect Fomu from
    // the host system.  Otherwise it would try to talk to
    // us over USB, which wouldn't work since we have no stack.
    assign usb_dp = 1'b0;
    assign usb_dn = 1'b0;
    assign usb_dp_pu = 1'b0;
    // Configure user pins so that we can detect the user connecting
    // 1-2 or 3-4 with conductive material.
    //
    // We do this by grounding user_2 and user_3, and configuring inputs
    // with pullups on user_1 and user_4.
    assign user_2 = 1'b0;
    assign user_3 = 1'b0;

    // Connect to system clock (with buffering)
    wire clk;
    SB_GB clk_gb (
        .USER_SIGNAL_TO_GLOBAL_BUFFER(clki),
        .GLOBAL_BUFFER_OUTPUT(clk)
    );

    // PyRTL module goes here:
    wire [3:0] colors;
    toplevel pyrtl_toplevel (
        .clk (clk),
        .in_1 (~user_1),
        .in_2 (~user_4),
        .red_o (colors[0]),
        .green_o (colors[1]),
        .blue_o (colors[2])
    );

    // Instantiate iCE40 LED driver hard logic, connecting up
    // counter state and LEDs.
    //
    // Note that it's possible to drive the LEDs directly,
    // however that is not current-limited and results in
    // overvolting the red LED.
    //
    // See also:
    // https://www.latticesemi.com/-/media/LatticeSemi/Documents/ApplicationNotes/IK/ICE40LEDDriverUsageGuide.ashx?document_id=50668
    SB_RGBA_DRV #(
        .CURRENT_MODE("0b1"),       // half current
        .RGB0_CURRENT("0b000011"),  // 4 mA
        .RGB1_CURRENT("0b000011"),  // 4 mA
        .RGB2_CURRENT("0b000011")   // 4 mA
    ) RGBA_DRIVER (
        .CURREN(1'b1),
        .RGBLEDEN(1'b1),
        .`REDPWM(colors[0]),      // Red
        .`GREENPWM(colors[1]),    // Green
        .`BLUEPWM(colors[2]),     // Blue
        .RGB0(rgb0),
        .RGB1(rgb1),
        .RGB2(rgb2)
    );

endmodule
// Generated automatically via PyRTL
// As one initial test of synthesis, map to FPGA with:
//   yosys -p "synth_xilinx -top toplevel" thisfile.v

module toplevel(clk, in_1, in_2, blue_o, green_o, red_o);
    input clk;
    input in_1;
    input in_2;
    output blue_o;
    output green_o;
    output red_o;

    reg[2:0] my_calculator_ctrl;
    reg[3:0] my_calculator_in_x;
    reg[3:0] my_calculator_in_y;
    reg[3:0] my_calculator_out_z;
    reg[26:0] tmp0;
    reg tmp5;
    reg tmp7;
    reg[15:0] tmp11;
    reg[15:0] tmp12;
    reg[15:0] tmp13;
    reg[15:0] tmp14;
    reg[15:0] tmp15;
    reg[15:0] tmp16;
    reg[15:0] tmp17;
    reg[15:0] tmp18;
    reg tmp19;
    reg[3:0] tmp8071;

    wire[15:0] _ver_out_tmp_0;
    wire[15:0] _ver_out_tmp_1;
    wire[15:0] _ver_out_tmp_2;
    wire[15:0] _ver_out_tmp_3;
    wire[15:0] _ver_out_tmp_4;
    wire[15:0] _ver_out_tmp_5;
    wire[15:0] _ver_out_tmp_6;
    wire[15:0] _ver_out_tmp_7;
    wire[15:0] _ver_out_tmp_8;
    wire[15:0] _ver_out_tmp_9;
    wire[15:0] _ver_out_tmp_10;
    wire[15:0] _ver_out_tmp_11;
    wire[15:0] _ver_out_tmp_12;
    wire[15:0] _ver_out_tmp_13;
    wire[15:0] _ver_out_tmp_14;
    wire[15:0] _ver_out_tmp_15;
    wire[15:0] _ver_out_tmp_16;
    wire[15:0] _ver_out_tmp_17;
    wire[15:0] _ver_out_tmp_18;
    wire[15:0] _ver_out_tmp_19;
    wire[15:0] _ver_out_tmp_20;
    wire[15:0] _ver_out_tmp_21;
    wire[15:0] _ver_out_tmp_22;
    wire[15:0] _ver_out_tmp_23;
    wire[15:0] _ver_out_tmp_24;
    wire[15:0] _ver_out_tmp_25;
    wire[15:0] _ver_out_tmp_26;
    wire[15:0] _ver_out_tmp_27;
    wire[15:0] _ver_out_tmp_28;
    wire[15:0] _ver_out_tmp_29;
    wire[15:0] _ver_out_tmp_30;
    wire[15:0] _ver_out_tmp_31;
    wire[15:0] _ver_out_tmp_32;
    wire[15:0] _ver_out_tmp_33;
    wire[15:0] _ver_out_tmp_34;
    wire[15:0] _ver_out_tmp_35;
    wire[15:0] _ver_out_tmp_36;
    wire[15:0] _ver_out_tmp_37;
    wire[15:0] _ver_out_tmp_38;
    wire[15:0] _ver_out_tmp_39;
    wire[15:0] _ver_out_tmp_40;
    wire[15:0] _ver_out_tmp_41;
    wire[15:0] _ver_out_tmp_42;
    wire[15:0] _ver_out_tmp_43;
    wire[15:0] _ver_out_tmp_44;
    wire[15:0] _ver_out_tmp_45;
    wire[15:0] _ver_out_tmp_46;
    wire[15:0] _ver_out_tmp_47;
    wire[15:0] _ver_out_tmp_48;
    wire[15:0] _ver_out_tmp_49;
    wire[15:0] _ver_out_tmp_50;
    wire[15:0] _ver_out_tmp_51;
    wire[15:0] _ver_out_tmp_52;
    wire[15:0] _ver_out_tmp_53;
    wire[15:0] _ver_out_tmp_54;
    wire[15:0] _ver_out_tmp_55;
    wire[15:0] _ver_out_tmp_56;
    wire[15:0] _ver_out_tmp_57;
    wire[15:0] _ver_out_tmp_58;
    wire[15:0] _ver_out_tmp_59;
    wire[15:0] _ver_out_tmp_60;
    wire[15:0] _ver_out_tmp_61;
    wire[15:0] _ver_out_tmp_62;
    wire[15:0] _ver_out_tmp_63;
    wire[15:0] _ver_out_tmp_64;
    wire[15:0] _ver_out_tmp_65;
    wire[15:0] _ver_out_tmp_66;
    wire[15:0] _ver_out_tmp_67;
    wire[15:0] _ver_out_tmp_68;
    wire[15:0] _ver_out_tmp_69;
    wire[15:0] _ver_out_tmp_70;
    wire[15:0] _ver_out_tmp_71;
    wire[15:0] _ver_out_tmp_72;
    wire[15:0] _ver_out_tmp_73;
    wire[15:0] _ver_out_tmp_74;
    wire[15:0] _ver_out_tmp_75;
    wire[15:0] _ver_out_tmp_76;
    wire[15:0] _ver_out_tmp_77;
    wire[15:0] _ver_out_tmp_78;
    wire[15:0] _ver_out_tmp_79;
    wire[15:0] _ver_out_tmp_80;
    wire[15:0] _ver_out_tmp_81;
    wire[15:0] _ver_out_tmp_82;
    wire[15:0] _ver_out_tmp_83;
    wire[15:0] _ver_out_tmp_84;
    wire[15:0] _ver_out_tmp_85;
    wire[15:0] _ver_out_tmp_86;
    wire[15:0] _ver_out_tmp_87;
    wire[15:0] _ver_out_tmp_88;
    wire[15:0] _ver_out_tmp_89;
    wire[15:0] _ver_out_tmp_90;
    wire[15:0] _ver_out_tmp_91;
    wire const_1_1;
    wire const_2_0;
    wire const_3_0;
    wire const_4_0;
    wire[2:0] const_5_4;
    wire[15:0] const_6_0;
    wire[15:0] const_7_2;
    wire[15:0] const_8_1;
    wire[15:0] const_9_0;
    wire[15:0] const_10_0;
    wire[15:0] const_11_0;
    wire[15:0] const_12_0;
    wire[15:0] const_13_1;
    wire const_14_0;
    wire const_15_1;
    wire const_16_0;
    wire[3:0] const_17_0;
    wire const_18_0;
    wire const_19_0;
    wire[3:0] const_20_15;
    wire const_21_1;
    wire const_22_0;
    wire[1:0] const_23_2;
    wire const_24_0;
    wire[1:0] const_25_3;
    wire const_26_0;
    wire const_27_0;
    wire const_28_0;
    wire const_29_0;
    wire const_30_0;
    wire const_31_0;
    wire[15:0] const_32_32767;
    wire const_34_0;
    wire const_35_0;
    wire const_36_0;
    wire const_37_0;
    wire const_38_0;
    wire[15:0] const_39_32767;
    wire const_41_0;
    wire const_42_0;
    wire const_43_0;
    wire const_44_0;
    wire const_45_0;
    wire[15:0] const_46_32767;
    wire const_48_0;
    wire const_49_0;
    wire const_50_0;
    wire const_51_0;
    wire const_52_0;
    wire[15:0] const_53_32767;
    wire[2:0] const_55_6;
    wire const_56_0;
    wire[2:0] const_57_7;
    wire const_58_0;
    wire[2:0] const_59_4;
    wire const_60_0;
    wire[2:0] const_61_5;
    wire const_62_0;
    wire const_63_0;
    wire const_64_0;
    wire const_65_0;
    wire const_66_0;
    wire const_67_0;
    wire const_68_0;
    wire[15:0] const_69_32767;
    wire const_71_0;
    wire const_72_0;
    wire const_73_0;
    wire const_74_0;
    wire const_75_0;
    wire const_76_0;
    wire[15:0] const_77_32767;
    wire const_79_0;
    wire const_80_0;
    wire const_81_0;
    wire const_82_0;
    wire const_83_0;
    wire const_84_0;
    wire[15:0] const_85_32767;
    wire const_87_0;
    wire const_88_0;
    wire const_89_0;
    wire const_90_0;
    wire const_91_0;
    wire const_92_0;
    wire[15:0] const_93_32767;
    wire[3:0] const_95_8;
    wire const_97_0;
    wire const_98_0;
    wire[14:0] const_99_32767;
    wire const_100_0;
    wire const_102_0;
    wire const_103_0;
    wire[14:0] const_104_32767;
    wire const_105_0;
    wire const_107_0;
    wire const_108_0;
    wire[14:0] const_109_32767;
    wire const_110_0;
    wire const_112_0;
    wire const_113_0;
    wire[14:0] const_114_32767;
    wire const_115_0;
    wire[1:0] const_116_2;
    wire const_117_0;
    wire[3:0] const_118_0;
    wire const_119_0;
    wire const_120_0;
    wire[3:0] const_121_15;
    wire const_122_1;
    wire const_123_0;
    wire[1:0] const_124_2;
    wire const_125_0;
    wire[1:0] const_126_3;
    wire const_127_0;
    wire const_128_0;
    wire const_129_0;
    wire const_130_0;
    wire const_131_0;
    wire const_132_0;
    wire[15:0] const_133_32767;
    wire const_135_0;
    wire const_136_0;
    wire const_137_0;
    wire const_138_0;
    wire const_139_0;
    wire[15:0] const_140_32767;
    wire const_142_0;
    wire const_143_0;
    wire const_144_0;
    wire const_145_0;
    wire const_146_0;
    wire[15:0] const_147_32767;
    wire const_149_0;
    wire const_150_0;
    wire const_151_0;
    wire const_152_0;
    wire const_153_0;
    wire[15:0] const_154_32767;
    wire[2:0] const_156_6;
    wire const_157_0;
    wire[2:0] const_158_7;
    wire const_159_0;
    wire[2:0] const_160_4;
    wire const_161_0;
    wire[2:0] const_162_5;
    wire const_163_0;
    wire const_164_0;
    wire const_165_0;
    wire const_166_0;
    wire const_167_0;
    wire const_168_0;
    wire const_169_0;
    wire[15:0] const_170_32767;
    wire const_172_0;
    wire const_173_0;
    wire const_174_0;
    wire const_175_0;
    wire const_176_0;
    wire const_177_0;
    wire[15:0] const_178_32767;
    wire const_180_0;
    wire const_181_0;
    wire const_182_0;
    wire const_183_0;
    wire const_184_0;
    wire const_185_0;
    wire[15:0] const_186_32767;
    wire const_188_0;
    wire const_189_0;
    wire const_190_0;
    wire const_191_0;
    wire const_192_0;
    wire const_193_0;
    wire[15:0] const_194_32767;
    wire[3:0] const_196_8;
    wire const_198_0;
    wire const_199_0;
    wire[14:0] const_200_32767;
    wire const_201_0;
    wire const_203_0;
    wire const_204_0;
    wire[14:0] const_205_32767;
    wire const_206_0;
    wire const_208_0;
    wire const_209_0;
    wire[14:0] const_210_32767;
    wire const_211_0;
    wire const_213_0;
    wire const_214_0;
    wire[14:0] const_215_32767;
    wire const_216_0;
    wire[1:0] const_217_3;
    wire const_218_0;
    wire const_219_0;
    wire const_220_0;
    wire const_221_0;
    wire const_222_0;
    wire const_223_0;
    wire const_224_0;
    wire const_225_0;
    wire const_226_0;
    wire const_227_0;
    wire const_228_0;
    wire const_229_0;
    wire const_230_0;
    wire const_231_0;
    wire const_232_0;
    wire const_233_0;
    wire const_234_0;
    wire const_235_0;
    wire const_236_0;
    wire const_237_0;
    wire const_238_0;
    wire const_239_0;
    wire const_240_0;
    wire const_242_0;
    wire const_243_0;
    wire[14:0] const_244_32767;
    wire const_245_0;
    wire const_247_0;
    wire const_248_0;
    wire[14:0] const_249_32767;
    wire const_250_0;
    wire const_252_0;
    wire const_253_0;
    wire[14:0] const_254_32767;
    wire const_255_0;
    wire const_257_0;
    wire const_258_0;
    wire[14:0] const_259_32767;
    wire const_260_0;
    wire const_262_0;
    wire const_263_0;
    wire[14:0] const_264_32767;
    wire const_265_0;
    wire const_267_0;
    wire const_268_0;
    wire[14:0] const_269_32767;
    wire const_270_0;
    wire const_272_0;
    wire const_273_0;
    wire[14:0] const_274_32767;
    wire const_275_0;
    wire const_277_0;
    wire const_278_0;
    wire[14:0] const_279_32767;
    wire const_280_0;
    wire const_281_0;
    wire const_282_0;
    wire const_283_0;
    wire const_284_0;
    wire const_285_0;
    wire const_286_0;
    wire const_287_0;
    wire const_288_0;
    wire const_289_0;
    wire const_290_0;
    wire[3:0] const_291_15;
    wire const_292_0;
    wire const_293_0;
    wire const_294_0;
    wire[3:0] const_295_8;
    wire const_296_0;
    wire const_298_0;
    wire const_299_0;
    wire[14:0] const_300_32767;
    wire const_301_0;
    wire const_303_0;
    wire const_304_0;
    wire[14:0] const_305_32767;
    wire const_306_0;
    wire const_308_0;
    wire const_309_0;
    wire[14:0] const_310_32767;
    wire const_311_0;
    wire const_313_0;
    wire const_314_0;
    wire[14:0] const_315_32767;
    wire const_316_0;
    wire[3:0] const_317_1;
    wire const_318_0;
    wire const_319_0;
    wire const_320_0;
    wire const_321_0;
    wire const_322_0;
    wire const_323_0;
    wire[15:0] const_324_32767;
    wire const_326_0;
    wire const_327_0;
    wire const_328_0;
    wire const_329_0;
    wire const_330_0;
    wire[15:0] const_331_32767;
    wire const_333_0;
    wire const_334_0;
    wire const_335_0;
    wire const_336_0;
    wire const_337_0;
    wire[15:0] const_338_32767;
    wire const_340_0;
    wire const_341_0;
    wire const_342_0;
    wire const_343_0;
    wire const_344_0;
    wire[15:0] const_345_32767;
    wire[3:0] const_347_4;
    wire const_348_0;
    wire const_350_0;
    wire const_351_0;
    wire[14:0] const_352_32767;
    wire const_353_0;
    wire const_354_0;
    wire const_355_0;
    wire const_356_0;
    wire const_357_0;
    wire const_358_0;
    wire const_359_0;
    wire[15:0] const_360_32767;
    wire const_363_0;
    wire const_364_0;
    wire[14:0] const_365_32767;
    wire const_366_0;
    wire const_367_0;
    wire const_368_0;
    wire const_369_0;
    wire const_370_0;
    wire const_371_0;
    wire const_372_0;
    wire[15:0] const_373_32767;
    wire const_376_0;
    wire const_377_0;
    wire[14:0] const_378_32767;
    wire const_379_0;
    wire const_380_0;
    wire const_381_0;
    wire const_382_0;
    wire const_383_0;
    wire const_384_0;
    wire const_385_0;
    wire[15:0] const_386_32767;
    wire const_389_0;
    wire const_390_0;
    wire[14:0] const_391_32767;
    wire const_392_0;
    wire const_393_0;
    wire const_394_0;
    wire const_395_0;
    wire const_396_0;
    wire const_397_0;
    wire const_398_0;
    wire[15:0] const_399_32767;
    wire[3:0] const_401_6;
    wire const_402_0;
    wire[1:0] const_403_0;
    wire const_404_0;
    wire const_405_0;
    wire const_406_0;
    wire const_407_0;
    wire[15:0] const_408_32767;
    wire[1:0] const_410_0;
    wire const_411_0;
    wire const_412_0;
    wire const_413_0;
    wire const_414_0;
    wire[15:0] const_415_32767;
    wire[1:0] const_417_0;
    wire const_418_0;
    wire const_419_0;
    wire const_420_0;
    wire const_421_0;
    wire[15:0] const_422_32767;
    wire[1:0] const_424_0;
    wire const_425_0;
    wire const_426_0;
    wire const_427_0;
    wire const_428_0;
    wire[15:0] const_429_32767;
    wire[3:0] const_431_2;
    wire const_432_0;
    wire const_433_0;
    wire const_434_0;
    wire const_435_0;
    wire const_436_0;
    wire const_437_0;
    wire[15:0] const_438_32767;
    wire const_440_0;
    wire const_441_0;
    wire const_442_0;
    wire const_443_0;
    wire const_444_0;
    wire[15:0] const_445_32767;
    wire const_447_0;
    wire const_448_0;
    wire const_449_0;
    wire const_450_0;
    wire const_451_0;
    wire[15:0] const_452_32767;
    wire const_454_0;
    wire const_455_0;
    wire const_456_0;
    wire const_457_0;
    wire const_458_0;
    wire[15:0] const_459_32767;
    wire const_461_0;
    wire const_462_0;
    wire const_463_0;
    wire const_464_0;
    wire const_465_0;
    wire[15:0] const_466_32767;
    wire const_468_0;
    wire const_469_0;
    wire const_470_0;
    wire const_471_0;
    wire const_472_0;
    wire[15:0] const_473_32767;
    wire const_475_0;
    wire const_476_0;
    wire const_477_0;
    wire const_478_0;
    wire const_479_0;
    wire[15:0] const_480_32767;
    wire const_482_0;
    wire const_483_0;
    wire const_484_0;
    wire const_485_0;
    wire const_486_0;
    wire[15:0] const_487_32767;
    wire const_489_0;
    wire const_490_0;
    wire const_491_0;
    wire const_492_0;
    wire const_493_0;
    wire[15:0] const_494_32767;
    wire const_496_0;
    wire const_497_0;
    wire const_498_0;
    wire const_499_0;
    wire const_500_0;
    wire[15:0] const_501_32767;
    wire const_503_0;
    wire const_504_0;
    wire const_505_0;
    wire const_506_0;
    wire const_507_0;
    wire[15:0] const_508_32767;
    wire const_510_0;
    wire const_511_0;
    wire const_512_0;
    wire const_513_0;
    wire const_514_0;
    wire[15:0] const_515_32767;
    wire[3:0] const_517_5;
    wire const_518_1;
    wire const_520_0;
    wire const_521_0;
    wire[14:0] const_522_32767;
    wire const_523_0;
    wire const_524_0;
    wire const_525_0;
    wire const_526_0;
    wire const_527_0;
    wire const_528_0;
    wire const_529_0;
    wire[15:0] const_530_32767;
    wire const_533_0;
    wire const_534_0;
    wire[14:0] const_535_32767;
    wire const_536_0;
    wire const_537_0;
    wire const_538_0;
    wire const_539_0;
    wire const_540_0;
    wire const_541_0;
    wire const_542_0;
    wire[15:0] const_543_32767;
    wire const_546_0;
    wire const_547_0;
    wire[14:0] const_548_32767;
    wire const_549_0;
    wire const_550_0;
    wire const_551_0;
    wire const_552_0;
    wire const_553_0;
    wire const_554_0;
    wire const_555_0;
    wire[15:0] const_556_32767;
    wire const_559_0;
    wire const_560_0;
    wire[14:0] const_561_32767;
    wire const_562_0;
    wire const_563_0;
    wire const_564_0;
    wire const_565_0;
    wire const_566_0;
    wire const_567_0;
    wire const_568_0;
    wire[15:0] const_569_32767;
    wire[3:0] const_571_0;
    wire const_572_0;
    wire[3:0] const_573_0;
    wire const_574_0;
    wire const_575_0;
    wire const_577_0;
    wire const_578_0;
    wire[14:0] const_579_32767;
    wire const_580_0;
    wire const_581_0;
    wire const_582_0;
    wire const_584_0;
    wire const_585_0;
    wire[14:0] const_586_32767;
    wire const_587_0;
    wire const_588_0;
    wire const_589_0;
    wire const_591_0;
    wire const_592_0;
    wire[14:0] const_593_32767;
    wire const_594_0;
    wire const_595_0;
    wire const_596_0;
    wire const_598_0;
    wire const_599_0;
    wire[14:0] const_600_32767;
    wire const_601_0;
    wire const_602_0;
    wire const_603_0;
    wire const_605_0;
    wire const_606_0;
    wire[14:0] const_607_32767;
    wire const_608_0;
    wire const_609_0;
    wire const_610_0;
    wire const_612_0;
    wire const_613_0;
    wire[14:0] const_614_32767;
    wire const_615_0;
    wire const_616_0;
    wire const_617_0;
    wire const_619_0;
    wire const_620_0;
    wire[14:0] const_621_32767;
    wire const_622_0;
    wire const_623_0;
    wire const_624_0;
    wire const_626_0;
    wire const_627_0;
    wire[14:0] const_628_32767;
    wire const_629_0;
    wire const_630_0;
    wire[3:0] const_631_6;
    wire const_632_1;
    wire const_633_0;
    wire const_635_0;
    wire const_636_0;
    wire[14:0] const_637_32767;
    wire const_638_0;
    wire const_639_0;
    wire const_640_0;
    wire const_642_0;
    wire const_643_0;
    wire[14:0] const_644_32767;
    wire const_645_0;
    wire const_646_0;
    wire const_647_0;
    wire const_649_0;
    wire const_650_0;
    wire[14:0] const_651_32767;
    wire const_652_0;
    wire const_653_0;
    wire const_654_0;
    wire const_656_0;
    wire const_657_0;
    wire[14:0] const_658_32767;
    wire const_659_0;
    wire const_660_0;
    wire const_661_0;
    wire const_663_0;
    wire const_664_0;
    wire[14:0] const_665_32767;
    wire const_666_0;
    wire const_667_0;
    wire const_668_0;
    wire const_670_0;
    wire const_671_0;
    wire[14:0] const_672_32767;
    wire const_673_0;
    wire const_674_0;
    wire const_675_0;
    wire const_677_0;
    wire const_678_0;
    wire[14:0] const_679_32767;
    wire const_680_0;
    wire const_681_0;
    wire const_682_0;
    wire const_684_0;
    wire const_685_0;
    wire[14:0] const_686_32767;
    wire const_687_0;
    wire const_688_0;
    wire[3:0] const_689_3;
    wire const_690_1;
    wire const_691_0;
    wire const_692_0;
    wire const_693_0;
    wire const_694_0;
    wire const_695_0;
    wire[15:0] const_696_32767;
    wire const_698_0;
    wire const_699_0;
    wire const_700_0;
    wire const_701_0;
    wire const_702_0;
    wire[15:0] const_703_32767;
    wire const_705_0;
    wire const_706_0;
    wire const_707_0;
    wire const_708_0;
    wire const_709_0;
    wire[15:0] const_710_32767;
    wire const_712_0;
    wire const_713_0;
    wire const_714_0;
    wire const_715_0;
    wire const_716_0;
    wire[15:0] const_717_32767;
    wire[3:0] const_719_0;
    wire[3:0] const_720_0;
    wire const_721_0;
    wire const_722_0;
    wire const_723_0;
    wire const_724_0;
    wire const_725_0;
    wire const_726_0;
    wire const_727_0;
    wire const_728_0;
    wire const_729_0;
    wire const_730_0;
    wire const_731_0;
    wire const_732_0;
    wire const_733_0;
    wire const_734_0;
    wire const_735_0;
    wire const_736_0;
    wire const_737_0;
    wire const_738_0;
    wire const_739_0;
    wire const_740_0;
    wire const_741_0;
    wire const_742_1;
    wire const_743_0;
    wire[1:0] const_744_2;
    wire const_745_0;
    wire[1:0] const_746_3;
    wire const_747_0;
    wire[3:0] const_748_15;
    wire[2:0] const_749_4;
    wire const_750_0;
    wire[2:0] const_751_5;
    wire const_752_0;
    wire[2:0] const_753_6;
    wire const_754_0;
    wire[2:0] const_755_7;
    wire const_756_0;
    wire[3:0] const_757_15;
    wire[3:0] const_758_8;
    wire[2:0] const_759_6;
    wire const_760_0;
    wire[2:0] const_761_7;
    wire const_762_0;
    wire[3:0] const_763_15;
    wire const_764_1;
    wire const_765_0;
    wire[2:0] const_766_2;
    wire[3:0] const_767_15;
    wire[1:0] const_768_2;
    wire const_769_0;
    wire[2:0] const_770_3;
    wire[1:0] const_771_3;
    wire const_772_0;
    wire[2:0] const_773_1;
    wire[3:0] const_774_15;
    wire[2:0] const_775_1;
    wire[3:0] const_776_15;
    wire const_781_0;
    wire const_782_0;
    wire const_783_0;
    wire const_784_0;
    wire[25:0] tmp1;
    wire[26:0] tmp2;
    wire[27:0] tmp3;
    wire[26:0] tmp4;
    wire tmp8;
    wire tmp10;
    wire tmp33;
    wire[2:0] tmp35;
    wire tmp36;
    wire tmp37;
    wire tmp73;
    wire[3:0] tmp90;
    wire tmp91;
    wire tmp92;
    wire tmp119;
    wire tmp131;
    wire tmp134;
    wire tmp135;
    wire tmp138;
    wire tmp139;
    wire[15:0] tmp141;
    wire[14:0] tmp143;
    wire tmp150;
    wire tmp152;
    wire[16:0] tmp158;
    wire tmp160;
    wire tmp161;
    wire tmp162;
    wire tmp166;
    wire[16:0] tmp183;
    wire tmp190;
    wire tmp192;
    wire tmp193;
    wire[15:0] tmp194;
    wire[15:0] tmp195;
    wire[14:0] tmp207;
    wire[15:0] tmp208;
    wire tmp217;
    wire[16:0] tmp225;
    wire tmp226;
    wire tmp228;
    wire tmp229;
    wire tmp232;
    wire tmp233;
    wire[16:0] tmp250;
    wire tmp251;
    wire tmp254;
    wire tmp255;
    wire tmp257;
    wire tmp258;
    wire tmp259;
    wire tmp260;
    wire[15:0] tmp261;
    wire[15:0] tmp262;
    wire tmp269;
    wire tmp273;
    wire[14:0] tmp274;
    wire[16:0] tmp292;
    wire tmp293;
    wire tmp318;
    wire tmp321;
    wire tmp325;
    wire[15:0] tmp329;
    wire[15:0] tmp342;
    wire tmp351;
    wire tmp354;
    wire[16:0] tmp359;
    wire tmp360;
    wire tmp362;
    wire tmp376;
    wire[16:0] tmp384;
    wire tmp385;
    wire tmp388;
    wire tmp389;
    wire tmp392;
    wire[15:0] tmp395;
    wire tmp410;
    wire tmp413;
    wire tmp414;
    wire tmp423;
    wire tmp424;
    wire tmp427;
    wire tmp459;
    wire[3:0] tmp520;
    wire tmp521;
    wire[3:0] tmp523;
    wire tmp524;
    wire tmp525;
    wire[17:0] tmp532;
    wire[16:0] tmp533;
    wire[15:0] tmp534;
    wire tmp558;
    wire tmp559;
    wire[16:0] tmp564;
    wire tmp565;
    wire tmp566;
    wire tmp568;
    wire tmp571;
    wire tmp573;
    wire tmp574;
    wire[16:0] tmp579;
    wire tmp586;
    wire tmp592;
    wire tmp593;
    wire tmp595;
    wire tmp599;
    wire[16:0] tmp604;
    wire tmp605;
    wire tmp608;
    wire tmp610;
    wire tmp611;
    wire tmp612;
    wire tmp613;
    wire tmp614;
    wire[15:0] tmp615;
    wire[15:0] tmp616;
    wire tmp642;
    wire tmp650;
    wire[17:0] tmp653;
    wire[16:0] tmp654;
    wire[15:0] tmp655;
    wire tmp667;
    wire tmp679;
    wire tmp680;
    wire[16:0] tmp685;
    wire tmp686;
    wire tmp689;
    wire tmp692;
    wire tmp693;
    wire tmp694;
    wire tmp695;
    wire tmp720;
    wire[16:0] tmp725;
    wire tmp726;
    wire tmp729;
    wire tmp730;
    wire tmp731;
    wire tmp732;
    wire tmp734;
    wire tmp735;
    wire[15:0] tmp736;
    wire[15:0] tmp737;
    wire tmp764;
    wire[16:0] tmp770;
    wire[17:0] tmp774;
    wire[16:0] tmp775;
    wire[15:0] tmp776;
    wire tmp782;
    wire tmp801;
    wire[16:0] tmp806;
    wire tmp807;
    wire tmp810;
    wire tmp813;
    wire tmp814;
    wire tmp815;
    wire tmp816;
    wire tmp834;
    wire tmp841;
    wire[16:0] tmp846;
    wire tmp847;
    wire tmp850;
    wire tmp851;
    wire tmp852;
    wire tmp853;
    wire tmp855;
    wire tmp856;
    wire[15:0] tmp857;
    wire[15:0] tmp858;
    wire tmp873;
    wire tmp889;
    wire[17:0] tmp895;
    wire[16:0] tmp896;
    wire[15:0] tmp897;
    wire tmp915;
    wire tmp918;
    wire tmp922;
    wire[16:0] tmp927;
    wire tmp928;
    wire tmp929;
    wire tmp930;
    wire tmp931;
    wire tmp934;
    wire tmp935;
    wire tmp936;
    wire tmp937;
    wire tmp943;
    wire tmp962;
    wire[16:0] tmp967;
    wire tmp968;
    wire tmp971;
    wire tmp974;
    wire tmp976;
    wire tmp977;
    wire[15:0] tmp978;
    wire[15:0] tmp979;
    wire tmp1010;
    wire tmp1051;
    wire tmp1057;
    wire tmp1083;
    wire tmp1086;
    wire[16:0] tmp1092;
    wire tmp1106;
    wire tmp1109;
    wire tmp1110;
    wire[2:0] tmp1112;
    wire tmp1113;
    wire tmp1132;
    wire tmp1133;
    wire tmp1141;
    wire tmp1166;
    wire[2:0] tmp1178;
    wire[3:0] tmp1179;
    wire tmp1180;
    wire tmp1183;
    wire tmp1184;
    wire tmp1187;
    wire tmp1188;
    wire[14:0] tmp1189;
    wire[16:0] tmp1195;
    wire tmp1196;
    wire tmp1202;
    wire tmp1208;
    wire tmp1214;
    wire tmp1221;
    wire tmp1233;
    wire tmp1236;
    wire tmp1240;
    wire[14:0] tmp1258;
    wire[15:0] tmp1259;
    wire tmp1265;
    wire tmp1268;
    wire[16:0] tmp1276;
    wire tmp1277;
    wire tmp1280;
    wire tmp1283;
    wire tmp1284;
    wire[16:0] tmp1301;
    wire tmp1302;
    wire tmp1305;
    wire tmp1306;
    wire tmp1307;
    wire tmp1308;
    wire tmp1309;
    wire tmp1310;
    wire tmp1311;
    wire[15:0] tmp1312;
    wire[15:0] tmp1313;
    wire[15:0] tmp1328;
    wire tmp1340;
    wire tmp1347;
    wire tmp1352;
    wire[16:0] tmp1370;
    wire tmp1377;
    wire tmp1379;
    wire tmp1380;
    wire[15:0] tmp1381;
    wire[15:0] tmp1397;
    wire tmp1403;
    wire[16:0] tmp1414;
    wire tmp1416;
    wire tmp1418;
    wire tmp1422;
    wire tmp1429;
    wire tmp1440;
    wire tmp1445;
    wire tmp1446;
    wire tmp1448;
    wire tmp1449;
    wire[15:0] tmp1451;
    wire tmp1464;
    wire tmp1467;
    wire tmp1470;
    wire tmp1471;
    wire tmp1484;
    wire tmp1542;
    wire tmp1555;
    wire tmp1561;
    wire tmp1594;
    wire tmp1597;
    wire tmp1598;
    wire[16:0] tmp1601;
    wire[16:0] tmp1604;
    wire[17:0] tmp1605;
    wire[16:0] tmp1606;
    wire[15:0] tmp1607;
    wire[16:0] tmp1624;
    wire tmp1625;
    wire tmp1629;
    wire tmp1632;
    wire[16:0] tmp1637;
    wire tmp1638;
    wire tmp1639;
    wire tmp1640;
    wire tmp1641;
    wire tmp1644;
    wire tmp1645;
    wire tmp1646;
    wire tmp1647;
    wire tmp1665;
    wire tmp1672;
    wire[16:0] tmp1677;
    wire tmp1678;
    wire tmp1681;
    wire tmp1684;
    wire tmp1686;
    wire tmp1687;
    wire[15:0] tmp1688;
    wire[15:0] tmp1689;
    wire tmp1701;
    wire[16:0] tmp1726;
    wire[16:0] tmp1729;
    wire[17:0] tmp1730;
    wire[16:0] tmp1731;
    wire[15:0] tmp1732;
    wire tmp1743;
    wire tmp1750;
    wire tmp1753;
    wire tmp1757;
    wire[16:0] tmp1762;
    wire tmp1763;
    wire tmp1764;
    wire tmp1765;
    wire tmp1766;
    wire tmp1769;
    wire tmp1770;
    wire tmp1771;
    wire tmp1772;
    wire[16:0] tmp1789;
    wire tmp1790;
    wire tmp1797;
    wire[16:0] tmp1802;
    wire tmp1803;
    wire tmp1806;
    wire tmp1809;
    wire tmp1811;
    wire tmp1812;
    wire[15:0] tmp1813;
    wire[15:0] tmp1814;
    wire tmp1841;
    wire tmp1846;
    wire tmp1849;
    wire[16:0] tmp1854;
    wire[17:0] tmp1855;
    wire[16:0] tmp1856;
    wire[15:0] tmp1857;
    wire tmp1866;
    wire tmp1882;
    wire[16:0] tmp1887;
    wire tmp1888;
    wire tmp1889;
    wire tmp1891;
    wire tmp1894;
    wire tmp1896;
    wire tmp1897;
    wire tmp1905;
    wire tmp1922;
    wire[16:0] tmp1927;
    wire tmp1928;
    wire tmp1931;
    wire tmp1933;
    wire tmp1934;
    wire tmp1935;
    wire tmp1936;
    wire tmp1937;
    wire[15:0] tmp1938;
    wire[15:0] tmp1939;
    wire[16:0] tmp1976;
    wire[16:0] tmp1979;
    wire[17:0] tmp1980;
    wire[16:0] tmp1981;
    wire[15:0] tmp1982;
    wire[16:0] tmp1999;
    wire tmp2006;
    wire tmp2007;
    wire[16:0] tmp2012;
    wire tmp2013;
    wire tmp2015;
    wire tmp2016;
    wire tmp2019;
    wire tmp2020;
    wire tmp2021;
    wire tmp2022;
    wire tmp2034;
    wire tmp2041;
    wire tmp2047;
    wire[16:0] tmp2052;
    wire tmp2053;
    wire tmp2056;
    wire tmp2057;
    wire tmp2059;
    wire tmp2061;
    wire tmp2062;
    wire[15:0] tmp2063;
    wire[15:0] tmp2064;
    wire tmp2078;
    wire tmp2081;
    wire tmp2099;
    wire tmp2100;
    wire[16:0] tmp2106;
    wire tmp2125;
    wire tmp2126;
    wire tmp2150;
    wire tmp2151;
    wire[2:0] tmp2209;
    wire tmp2235;
    wire[16:0] tmp2240;
    wire tmp2247;
    wire tmp2260;
    wire tmp2261;
    wire tmp2281;
    wire tmp2286;
    wire tmp2287;
    wire tmp2322;
    wire tmp2343;
    wire tmp2347;
    wire tmp2348;
    wire[16:0] tmp2353;
    wire[16:0] tmp2365;
    wire tmp2366;
    wire tmp2369;
    wire tmp2373;
    wire tmp2374;
    wire tmp2387;
    wire tmp2390;
    wire tmp2391;
    wire tmp2395;
    wire tmp2398;
    wire tmp2399;
    wire tmp2410;
    wire tmp2411;
    wire tmp2412;
    wire tmp2423;
    wire tmp2424;
    wire tmp2425;
    wire tmp2426;
    wire tmp2427;
    wire tmp2428;
    wire tmp2429;
    wire tmp2430;
    wire tmp2453;
    wire[16:0] tmp2458;
    wire tmp2466;
    wire[15:0] tmp2474;
    wire tmp2486;
    wire[16:0] tmp2492;
    wire[15:0] tmp2512;
    wire tmp2524;
    wire[16:0] tmp2527;
    wire[16:0] tmp2530;
    wire[15:0] tmp2531;
    wire[16:0] tmp2549;
    wire[15:0] tmp2550;
    wire tmp2561;
    wire[16:0] tmp2565;
    wire[15:0] tmp2569;
    wire tmp2581;
    wire[15:0] tmp2588;
    wire[16:0] tmp2606;
    wire[15:0] tmp2607;
    wire tmp2610;
    wire tmp2625;
    wire tmp2627;
    wire tmp2643;
    wire tmp2644;
    wire tmp2645;
    wire tmp2646;
    wire tmp2649;
    wire tmp2681;
    wire tmp2722;
    wire tmp2736;
    wire tmp2747;
    wire tmp2756;
    wire tmp2759;
    wire tmp2760;
    wire tmp2764;
    wire tmp2775;
    wire tmp2807;
    wire tmp2811;
    wire tmp2812;
    wire tmp2826;
    wire[15:0] tmp2870;
    wire tmp2885;
    wire[15:0] tmp2887;
    wire[16:0] tmp2935;
    wire tmp2936;
    wire tmp2937;
    wire tmp2939;
    wire tmp2942;
    wire tmp2943;
    wire tmp2944;
    wire[15:0] tmp2948;
    wire[16:0] tmp2951;
    wire tmp2952;
    wire tmp2953;
    wire tmp2954;
    wire tmp2955;
    wire tmp2958;
    wire tmp2959;
    wire tmp2960;
    wire tmp2961;
    wire[16:0] tmp2968;
    wire tmp2969;
    wire tmp2970;
    wire tmp2972;
    wire tmp2975;
    wire tmp2976;
    wire tmp2977;
    wire tmp2978;
    wire[15:0] tmp2982;
    wire[16:0] tmp2985;
    wire tmp2986;
    wire tmp2987;
    wire tmp2988;
    wire tmp2989;
    wire tmp2992;
    wire tmp2993;
    wire tmp2994;
    wire tmp2995;
    wire tmp3029;
    wire tmp3145;
    wire tmp3196;
    wire tmp3215;
    wire[15:0] tmp3253;
    wire tmp3263;
    wire[16:0] tmp3270;
    wire tmp3271;
    wire tmp3274;
    wire tmp3278;
    wire tmp3284;
    wire tmp3287;
    wire tmp3290;
    wire[15:0] tmp3307;
    wire[15:0] tmp3327;
    wire tmp3345;
    wire tmp3347;
    wire tmp3348;
    wire tmp3351;
    wire tmp3360;
    wire tmp3361;
    wire tmp3373;
    wire tmp3376;
    wire tmp3379;
    wire tmp3397;
    wire tmp3413;
    wire tmp3419;
    wire tmp3435;
    wire tmp3453;
    wire[16:0] tmp3480;
    wire tmp3486;
    wire tmp3496;
    wire tmp3506;
    wire tmp3521;
    wire tmp3526;
    wire[15:0] tmp3528;
    wire[16:0] tmp3550;
    wire tmp3553;
    wire tmp3554;
    wire tmp3557;
    wire tmp3558;
    wire tmp3559;
    wire tmp3566;
    wire tmp3569;
    wire tmp3570;
    wire tmp3571;
    wire tmp3572;
    wire[16:0] tmp3575;
    wire tmp3576;
    wire tmp3579;
    wire tmp3582;
    wire tmp3583;
    wire tmp3584;
    wire tmp3585;
    wire[16:0] tmp3588;
    wire tmp3589;
    wire tmp3592;
    wire tmp3595;
    wire tmp3596;
    wire tmp3597;
    wire tmp3598;
    wire[14:0] tmp3599;
    wire[15:0] tmp3602;
    wire[16:0] tmp3605;
    wire tmp3606;
    wire tmp3608;
    wire tmp3609;
    wire tmp3612;
    wire tmp3613;
    wire[14:0] tmp3614;
    wire[16:0] tmp3620;
    wire tmp3621;
    wire tmp3624;
    wire tmp3627;
    wire tmp3628;
    wire tmp3630;
    wire[16:0] tmp3635;
    wire tmp3636;
    wire tmp3638;
    wire tmp3639;
    wire tmp3640;
    wire tmp3642;
    wire tmp3643;
    wire[16:0] tmp3650;
    wire tmp3651;
    wire tmp3654;
    wire tmp3657;
    wire tmp3658;
    wire tmp3694;
    wire tmp3713;
    wire[16:0] tmp3719;
    wire[1:0] tmp3721;
    wire[17:0] tmp3722;
    wire[17:0] tmp3725;
    wire[18:0] tmp3726;
    wire[17:0] tmp3727;
    wire[15:0] tmp3728;
    wire[16:0] tmp3733;
    wire tmp3734;
    wire tmp3737;
    wire[15:0] tmp3742;
    wire[17:0] tmp3745;
    wire tmp3746;
    wire tmp3752;
    wire tmp3753;
    wire[16:0] tmp3758;
    wire tmp3759;
    wire tmp3760;
    wire tmp3762;
    wire tmp3765;
    wire tmp3766;
    wire[16:0] tmp3773;
    wire tmp3777;
    wire tmp3780;
    wire[17:0] tmp3785;
    wire tmp3786;
    wire tmp3788;
    wire tmp3793;
    wire[16:0] tmp3798;
    wire tmp3802;
    wire[15:0] tmp3810;
    wire[17:0] tmp3856;
    wire[18:0] tmp3860;
    wire[17:0] tmp3861;
    wire[16:0] tmp3867;
    wire tmp3880;
    wire[16:0] tmp3892;
    wire tmp3893;
    wire tmp3901;
    wire[17:0] tmp3919;
    wire tmp3921;
    wire tmp3922;
    wire tmp3926;
    wire tmp3937;
    wire tmp3939;
    wire tmp3940;
    wire tmp3941;
    wire[15:0] tmp3943;
    wire[15:0] tmp3944;
    wire[16:0] tmp3987;
    wire tmp3988;
    wire[17:0] tmp3990;
    wire tmp3991;
    wire[17:0] tmp3995;
    wire[15:0] tmp3996;
    wire[16:0] tmp4001;
    wire tmp4008;
    wire[17:0] tmp4013;
    wire tmp4014;
    wire tmp4016;
    wire tmp4017;
    wire tmp4021;
    wire[16:0] tmp4026;
    wire tmp4027;
    wire tmp4030;
    wire tmp4033;
    wire tmp4035;
    wire tmp4036;
    wire[16:0] tmp4041;
    wire tmp4045;
    wire[17:0] tmp4053;
    wire tmp4054;
    wire tmp4056;
    wire tmp4057;
    wire tmp4060;
    wire tmp4061;
    wire[16:0] tmp4066;
    wire tmp4067;
    wire tmp4070;
    wire tmp4071;
    wire tmp4072;
    wire tmp4073;
    wire tmp4076;
    wire[15:0] tmp4077;
    wire[15:0] tmp4078;
    wire[1:0] tmp4123;
    wire[17:0] tmp4127;
    wire[18:0] tmp4128;
    wire[17:0] tmp4129;
    wire[15:0] tmp4130;
    wire[16:0] tmp4135;
    wire tmp4142;
    wire tmp4153;
    wire tmp4155;
    wire tmp4168;
    wire tmp4169;
    wire tmp4170;
    wire tmp4182;
    wire[17:0] tmp4187;
    wire tmp4207;
    wire tmp4209;
    wire tmp4210;
    wire[15:0] tmp4212;
    wire[16:0] tmp4233;
    wire tmp4234;
    wire tmp4237;
    wire tmp4240;
    wire[16:0] tmp4243;
    wire tmp4244;
    wire tmp4247;
    wire tmp4250;
    wire tmp4251;
    wire[16:0] tmp4254;
    wire tmp4255;
    wire tmp4257;
    wire tmp4258;
    wire tmp4261;
    wire tmp4262;
    wire[16:0] tmp4265;
    wire tmp4266;
    wire tmp4269;
    wire tmp4272;
    wire tmp4273;
    wire tmp4395;
    wire tmp4413;
    wire tmp4469;
    wire tmp4477;
    wire tmp4480;
    wire tmp4481;
    wire tmp4483;
    wire[13:0] tmp4484;
    wire[15:0] tmp4485;
    wire tmp4494;
    wire tmp4497;
    wire[16:0] tmp4502;
    wire tmp4503;
    wire tmp4504;
    wire tmp4505;
    wire tmp4506;
    wire tmp4509;
    wire tmp4510;
    wire[16:0] tmp4527;
    wire tmp4528;
    wire tmp4531;
    wire tmp4534;
    wire tmp4535;
    wire tmp4536;
    wire tmp4537;
    wire[15:0] tmp4538;
    wire[15:0] tmp4539;
    wire[16:0] tmp4542;
    wire tmp4543;
    wire tmp4546;
    wire tmp4547;
    wire tmp4548;
    wire tmp4549;
    wire tmp4550;
    wire[16:0] tmp4553;
    wire tmp4554;
    wire tmp4557;
    wire tmp4560;
    wire tmp4561;
    wire[13:0] tmp4562;
    wire[15:0] tmp4563;
    wire tmp4573;
    wire tmp4575;
    wire[16:0] tmp4580;
    wire tmp4581;
    wire tmp4582;
    wire tmp4583;
    wire tmp4584;
    wire tmp4587;
    wire tmp4588;
    wire tmp4594;
    wire[16:0] tmp4605;
    wire tmp4606;
    wire tmp4609;
    wire tmp4612;
    wire tmp4613;
    wire tmp4614;
    wire tmp4615;
    wire[15:0] tmp4616;
    wire[15:0] tmp4617;
    wire[16:0] tmp4620;
    wire tmp4621;
    wire tmp4623;
    wire tmp4624;
    wire tmp4625;
    wire tmp4626;
    wire tmp4627;
    wire tmp4628;
    wire tmp4635;
    wire tmp4638;
    wire tmp4639;
    wire[13:0] tmp4640;
    wire[15:0] tmp4641;
    wire tmp4652;
    wire[16:0] tmp4658;
    wire tmp4659;
    wire tmp4660;
    wire tmp4661;
    wire tmp4662;
    wire tmp4665;
    wire tmp4666;
    wire[16:0] tmp4683;
    wire tmp4684;
    wire tmp4687;
    wire tmp4690;
    wire tmp4691;
    wire tmp4692;
    wire tmp4693;
    wire[15:0] tmp4694;
    wire[15:0] tmp4695;
    wire[16:0] tmp4698;
    wire tmp4699;
    wire tmp4702;
    wire tmp4703;
    wire tmp4704;
    wire tmp4705;
    wire tmp4706;
    wire tmp4713;
    wire tmp4716;
    wire tmp4717;
    wire[13:0] tmp4718;
    wire[15:0] tmp4719;
    wire tmp4725;
    wire tmp4729;
    wire[16:0] tmp4736;
    wire tmp4737;
    wire tmp4740;
    wire tmp4743;
    wire tmp4744;
    wire[16:0] tmp4761;
    wire tmp4762;
    wire tmp4765;
    wire tmp4766;
    wire tmp4767;
    wire tmp4768;
    wire tmp4769;
    wire tmp4770;
    wire tmp4771;
    wire[15:0] tmp4772;
    wire[15:0] tmp4773;
    wire[16:0] tmp4776;
    wire tmp4777;
    wire tmp4780;
    wire tmp4781;
    wire tmp4782;
    wire tmp4783;
    wire tmp4784;
    wire tmp4860;
    wire tmp4886;
    wire[14:0] tmp4887;
    wire[15:0] tmp4890;
    wire[14:0] tmp4915;
    wire tmp4916;
    wire tmp4971;
    wire tmp4999;
    wire tmp5011;
    wire tmp5013;
    wire tmp5102;
    wire[14:0] tmp5139;
    wire[16:0] tmp5145;
    wire tmp5146;
    wire tmp5164;
    wire[16:0] tmp5170;
    wire tmp5173;
    wire[16:0] tmp5182;
    wire tmp5187;
    wire tmp5189;
    wire tmp5192;
    wire[15:0] tmp5193;
    wire tmp5209;
    wire tmp5219;
    wire tmp5271;
    wire tmp5272;
    wire[15:0] tmp5274;
    wire[14:0] tmp5301;
    wire tmp5311;
    wire tmp5323;
    wire tmp5326;
    wire tmp5327;
    wire tmp5345;
    wire tmp5352;
    wire tmp5353;
    wire[15:0] tmp5356;
    wire tmp5395;
    wire[16:0] tmp5400;
    wire tmp5401;
    wire tmp5402;
    wire tmp5417;
    wire tmp5420;
    wire[16:0] tmp5425;
    wire tmp5426;
    wire tmp5432;
    wire tmp5435;
    wire[14:0] tmp5463;
    wire[15:0] tmp5464;
    wire[16:0] tmp5481;
    wire tmp5482;
    wire tmp5483;
    wire tmp5484;
    wire tmp5485;
    wire tmp5488;
    wire tmp5489;
    wire tmp5495;
    wire[16:0] tmp5506;
    wire tmp5507;
    wire tmp5508;
    wire tmp5510;
    wire tmp5513;
    wire tmp5514;
    wire tmp5515;
    wire tmp5516;
    wire[15:0] tmp5517;
    wire[15:0] tmp5518;
    wire[16:0] tmp5521;
    wire tmp5522;
    wire tmp5525;
    wire tmp5526;
    wire tmp5527;
    wire tmp5528;
    wire tmp5550;
    wire tmp5573;
    wire tmp5576;
    wire tmp5580;
    wire tmp5581;
    wire[16:0] tmp5587;
    wire tmp5588;
    wire tmp5591;
    wire tmp5592;
    wire tmp5593;
    wire tmp5594;
    wire tmp5595;
    wire[14:0] tmp5596;
    wire[15:0] tmp5597;
    wire tmp5603;
    wire tmp5606;
    wire tmp5607;
    wire tmp5609;
    wire[16:0] tmp5614;
    wire tmp5615;
    wire tmp5616;
    wire tmp5617;
    wire tmp5618;
    wire tmp5621;
    wire tmp5622;
    wire[16:0] tmp5627;
    wire tmp5628;
    wire tmp5631;
    wire tmp5634;
    wire[16:0] tmp5639;
    wire tmp5640;
    wire tmp5643;
    wire tmp5646;
    wire tmp5647;
    wire tmp5648;
    wire tmp5649;
    wire[15:0] tmp5650;
    wire[15:0] tmp5651;
    wire[16:0] tmp5654;
    wire tmp5655;
    wire tmp5658;
    wire tmp5659;
    wire tmp5660;
    wire tmp5661;
    wire tmp5662;
    wire[14:0] tmp5663;
    wire[16:0] tmp5669;
    wire tmp5670;
    wire tmp5673;
    wire[16:0] tmp5681;
    wire tmp5683;
    wire tmp5689;
    wire[16:0] tmp5694;
    wire tmp5701;
    wire[16:0] tmp5706;
    wire tmp5707;
    wire[15:0] tmp5718;
    wire[16:0] tmp5721;
    wire tmp5722;
    wire tmp5725;
    wire tmp5726;
    wire tmp5727;
    wire tmp5728;
    wire tmp5729;
    wire[14:0] tmp5730;
    wire[15:0] tmp5731;
    wire tmp5740;
    wire[16:0] tmp5748;
    wire tmp5749;
    wire tmp5752;
    wire tmp5755;
    wire tmp5756;
    wire tmp5768;
    wire[16:0] tmp5773;
    wire tmp5774;
    wire tmp5777;
    wire tmp5778;
    wire tmp5779;
    wire tmp5780;
    wire tmp5781;
    wire tmp5782;
    wire tmp5783;
    wire[15:0] tmp5784;
    wire[15:0] tmp5785;
    wire[16:0] tmp5788;
    wire tmp5789;
    wire tmp5792;
    wire tmp5793;
    wire tmp5794;
    wire tmp5795;
    wire tmp5796;
    wire[15:0] tmp5798;
    wire[16:0] tmp5803;
    wire tmp5804;
    wire[16:0] tmp5815;
    wire tmp5817;
    wire[16:0] tmp5828;
    wire tmp5829;
    wire tmp5835;
    wire[16:0] tmp5840;
    wire tmp5844;
    wire tmp5846;
    wire tmp5847;
    wire[15:0] tmp5851;
    wire[16:0] tmp5855;
    wire tmp5856;
    wire tmp5859;
    wire tmp5860;
    wire tmp5861;
    wire tmp5862;
    wire tmp5863;
    wire[14:0] tmp5864;
    wire[15:0] tmp5865;
    wire tmp5871;
    wire tmp5874;
    wire[16:0] tmp5882;
    wire tmp5883;
    wire tmp5886;
    wire tmp5889;
    wire tmp5890;
    wire tmp5899;
    wire[16:0] tmp5907;
    wire tmp5908;
    wire tmp5911;
    wire tmp5912;
    wire tmp5913;
    wire tmp5914;
    wire tmp5915;
    wire tmp5916;
    wire tmp5917;
    wire[15:0] tmp5918;
    wire[15:0] tmp5919;
    wire[16:0] tmp5922;
    wire tmp5923;
    wire tmp5926;
    wire tmp5927;
    wire tmp5928;
    wire tmp5929;
    wire tmp5930;
    wire[14:0] tmp5931;
    wire[15:0] tmp5932;
    wire tmp5941;
    wire tmp5952;
    wire tmp5956;
    wire tmp5957;
    wire[16:0] tmp5962;
    wire tmp5982;
    wire[15:0] tmp5986;
    wire[16:0] tmp5989;
    wire tmp5990;
    wire tmp5993;
    wire tmp5994;
    wire tmp5995;
    wire tmp5996;
    wire tmp5997;
    wire tmp6072;
    wire tmp6083;
    wire tmp6100;
    wire tmp6107;
    wire tmp6109;
    wire tmp6127;
    wire tmp6128;
    wire tmp6149;
    wire tmp6152;
    wire tmp6159;
    wire tmp6164;
    wire tmp6165;
    wire tmp6167;
    wire tmp6168;
    wire[15:0] tmp6169;
    wire tmp6183;
    wire tmp6221;
    wire[16:0] tmp6227;
    wire[1:0] tmp6229;
    wire[17:0] tmp6233;
    wire[15:0] tmp6236;
    wire[17:0] tmp6253;
    wire tmp6257;
    wire tmp6260;
    wire tmp6261;
    wire tmp6270;
    wire tmp6273;
    wire tmp6276;
    wire tmp6294;
    wire tmp6297;
    wire tmp6301;
    wire[16:0] tmp6306;
    wire tmp6307;
    wire tmp6310;
    wire tmp6312;
    wire tmp6316;
    wire tmp6366;
    wire tmp6367;
    wire tmp6369;
    wire[1:0] tmp6377;
    wire[17:0] tmp6381;
    wire[18:0] tmp6382;
    wire tmp6390;
    wire tmp6408;
    wire tmp6430;
    wire[16:0] tmp6440;
    wire tmp6462;
    wire tmp6463;
    wire tmp6517;
    wire[16:0] tmp6523;
    wire[17:0] tmp6526;
    wire tmp6542;
    wire tmp6543;
    wire[17:0] tmp6549;
    wire tmp6550;
    wire tmp6553;
    wire tmp6556;
    wire[16:0] tmp6562;
    wire tmp6563;
    wire tmp6566;
    wire tmp6569;
    wire[16:0] tmp6577;
    wire tmp6578;
    wire tmp6590;
    wire tmp6591;
    wire tmp6593;
    wire tmp6596;
    wire tmp6597;
    wire[16:0] tmp6602;
    wire tmp6603;
    wire tmp6605;
    wire tmp6606;
    wire tmp6607;
    wire tmp6608;
    wire[15:0] tmp6613;
    wire tmp6633;
    wire tmp6634;
    wire tmp6656;
    wire tmp6657;
    wire tmp6665;
    wire tmp6690;
    wire[16:0] tmp6758;
    wire[16:0] tmp6759;
    wire tmp6765;
    wire tmp6772;
    wire[16:0] tmp6781;
    wire[17:0] tmp6784;
    wire tmp6785;
    wire tmp6786;
    wire tmp6787;
    wire tmp6788;
    wire tmp6791;
    wire[1:0] tmp6808;
    wire[16:0] tmp6813;
    wire tmp6825;
    wire[16:0] tmp6834;
    wire[17:0] tmp6838;
    wire tmp6839;
    wire tmp6840;
    wire tmp6841;
    wire tmp6842;
    wire tmp6843;
    wire tmp6844;
    wire tmp6845;
    wire tmp6846;
    wire[16:0] tmp6851;
    wire[16:0] tmp6864;
    wire[16:0] tmp6865;
    wire[16:0] tmp6887;
    wire[16:0] tmp6889;
    wire[16:0] tmp6890;
    wire[17:0] tmp6893;
    wire tmp6894;
    wire tmp6895;
    wire tmp6896;
    wire tmp6897;
    wire tmp6900;
    wire tmp6901;
    wire tmp6910;
    wire tmp6913;
    wire tmp6931;
    wire tmp6935;
    wire tmp6936;
    wire[16:0] tmp6945;
    wire[17:0] tmp6948;
    wire tmp6949;
    wire tmp6950;
    wire tmp6951;
    wire tmp6952;
    wire tmp6953;
    wire tmp6954;
    wire tmp6955;
    wire tmp6956;
    wire tmp7020;
    wire tmp7031;
    wire[15:0] tmp7139;
    wire tmp7140;
    wire[16:0] tmp7142;
    wire tmp7154;
    wire[16:0] tmp7163;
    wire[17:0] tmp7167;
    wire tmp7168;
    wire tmp7169;
    wire tmp7170;
    wire tmp7171;
    wire tmp7172;
    wire tmp7173;
    wire tmp7174;
    wire tmp7175;
    wire tmp7176;
    wire tmp7177;
    wire tmp7185;
    wire tmp7186;
    wire[16:0] tmp7198;
    wire[15:0] tmp7200;
    wire tmp7201;
    wire[16:0] tmp7203;
    wire[16:0] tmp7225;
    wire[17:0] tmp7228;
    wire tmp7229;
    wire tmp7230;
    wire tmp7231;
    wire tmp7232;
    wire tmp7235;
    wire tmp7236;
    wire tmp7237;
    wire tmp7238;
    wire tmp7250;
    wire[16:0] tmp7254;
    wire[16:0] tmp7259;
    wire[16:0] tmp7260;
    wire[15:0] tmp7261;
    wire tmp7262;
    wire[16:0] tmp7264;
    wire[16:0] tmp7280;
    wire[17:0] tmp7289;
    wire tmp7290;
    wire tmp7291;
    wire tmp7292;
    wire tmp7293;
    wire tmp7294;
    wire tmp7295;
    wire tmp7296;
    wire tmp7297;
    wire tmp7298;
    wire tmp7299;
    wire[16:0] tmp7320;
    wire[16:0] tmp7321;
    wire[15:0] tmp7322;
    wire tmp7323;
    wire[16:0] tmp7325;
    wire[16:0] tmp7346;
    wire[17:0] tmp7350;
    wire tmp7351;
    wire tmp7352;
    wire tmp7353;
    wire tmp7354;
    wire tmp7357;
    wire tmp7358;
    wire tmp7359;
    wire tmp7360;
    wire[14:0] tmp7397;
    wire tmp7398;
    wire[15:0] tmp7400;
    wire tmp7419;
    wire[14:0] tmp7420;
    wire tmp7421;
    wire[15:0] tmp7423;
    wire tmp7435;
    wire[14:0] tmp7443;
    wire tmp7444;
    wire[15:0] tmp7446;
    wire[14:0] tmp7466;
    wire tmp7467;
    wire[15:0] tmp7469;
    wire[16:0] tmp7495;
    wire tmp7511;
    wire tmp7515;
    wire tmp7538;
    wire tmp7558;
    wire tmp7564;
    wire[14:0] tmp7565;
    wire tmp7572;
    wire tmp7577;
    wire tmp7587;
    wire tmp7590;
    wire tmp7591;
    wire[16:0] tmp7596;
    wire tmp7615;
    wire tmp7617;
    wire tmp7618;
    wire[15:0] tmp7620;
    wire tmp7628;
    wire[14:0] tmp7641;
    wire tmp7651;
    wire tmp7654;
    wire tmp7660;
    wire tmp7666;
    wire tmp7675;
    wire[16:0] tmp7684;
    wire tmp7688;
    wire tmp7692;
    wire[15:0] tmp7695;
    wire[14:0] tmp7717;
    wire[15:0] tmp7718;
    wire[16:0] tmp7735;
    wire tmp7736;
    wire tmp7738;
    wire tmp7739;
    wire tmp7742;
    wire tmp7743;
    wire[16:0] tmp7760;
    wire tmp7761;
    wire tmp7764;
    wire tmp7765;
    wire tmp7767;
    wire tmp7768;
    wire tmp7769;
    wire tmp7770;
    wire[15:0] tmp7771;
    wire[15:0] tmp7772;
    wire tmp7785;
    wire tmp7790;
    wire tmp7809;
    wire tmp7810;
    wire tmp7818;
    wire tmp7827;
    wire tmp7830;
    wire[15:0] tmp7863;
    wire[15:0] tmp7864;
    wire[15:0] tmp7865;
    wire[15:0] tmp7866;
    wire[15:0] tmp7867;
    wire[15:0] tmp7868;
    wire[15:0] tmp7869;
    wire[15:0] tmp7870;
    wire[15:0] tmp7871;
    wire[15:0] tmp7872;
    wire[15:0] tmp7873;
    wire[15:0] tmp7874;
    wire[15:0] tmp7875;
    wire[15:0] tmp7876;
    wire[15:0] tmp7877;
    wire[15:0] tmp7878;
    wire[15:0] tmp7879;
    wire[15:0] tmp7880;
    wire[15:0] tmp7881;
    wire[15:0] tmp7882;
    wire[15:0] tmp7883;
    wire[15:0] tmp7884;
    wire[15:0] tmp7885;
    wire[15:0] tmp7886;
    wire[15:0] tmp7887;
    wire[15:0] tmp7888;
    wire[15:0] tmp7889;
    wire[15:0] tmp7890;
    wire[15:0] tmp7891;
    wire[15:0] tmp7892;
    wire[15:0] tmp7893;
    wire[15:0] tmp7894;
    wire[15:0] tmp7895;
    wire[15:0] tmp7896;
    wire[15:0] tmp7897;
    wire[15:0] tmp7898;
    wire[15:0] tmp7899;
    wire[15:0] tmp7900;
    wire[15:0] tmp7901;
    wire[15:0] tmp7902;
    wire[15:0] tmp7903;
    wire[15:0] tmp7904;
    wire[15:0] tmp7905;
    wire[15:0] tmp7906;
    wire[15:0] tmp7907;
    wire[15:0] tmp7908;
    wire[15:0] tmp7909;
    wire[15:0] tmp7910;
    wire[15:0] tmp7911;
    wire[15:0] tmp7912;
    wire[15:0] tmp7913;
    wire[15:0] tmp7914;
    wire[15:0] tmp7915;
    wire[15:0] tmp7916;
    wire[15:0] tmp7917;
    wire[15:0] tmp7918;
    wire[15:0] tmp7919;
    wire[15:0] tmp7920;
    wire[15:0] tmp7921;
    wire[15:0] tmp7922;
    wire[15:0] tmp7923;
    wire[15:0] tmp7924;
    wire[15:0] tmp7925;
    wire[15:0] tmp7926;
    wire[15:0] tmp7927;
    wire[15:0] tmp7928;
    wire[15:0] tmp7929;
    wire[15:0] tmp7930;
    wire[15:0] tmp7931;
    wire[15:0] tmp7932;
    wire[15:0] tmp7933;
    wire[15:0] tmp7934;
    wire[15:0] tmp7935;
    wire[15:0] tmp7936;
    wire[15:0] tmp7937;
    wire[15:0] tmp7938;
    wire[15:0] tmp7939;
    wire[15:0] tmp7940;
    wire[15:0] tmp7941;
    wire[15:0] tmp7942;
    wire[15:0] tmp7943;
    wire[15:0] tmp7944;
    wire[15:0] tmp7945;
    wire[15:0] tmp7946;
    wire[15:0] tmp7947;
    wire[15:0] tmp7948;
    wire[15:0] tmp7949;
    wire[15:0] tmp7950;
    wire[15:0] tmp7951;
    wire[15:0] tmp7952;
    wire[15:0] tmp7953;
    wire[15:0] tmp7954;
    wire[15:0] tmp7955;
    wire[15:0] tmp7956;
    wire[15:0] tmp7957;
    wire[15:0] tmp7958;
    wire[15:0] tmp7959;
    wire[15:0] tmp7960;
    wire[15:0] tmp7961;
    wire[15:0] tmp7962;
    wire[15:0] tmp7963;
    wire[15:0] tmp7964;
    wire[15:0] tmp7965;
    wire[15:0] tmp7966;
    wire[15:0] tmp7967;
    wire[15:0] tmp7968;
    wire[15:0] tmp7969;
    wire[15:0] tmp7970;
    wire[15:0] tmp7971;
    wire[15:0] tmp7972;
    wire[15:0] tmp7973;
    wire[15:0] tmp7974;
    wire[15:0] tmp7975;
    wire[15:0] tmp7976;
    wire[15:0] tmp7977;
    wire[15:0] tmp7978;
    wire[15:0] tmp7979;
    wire[15:0] tmp7980;
    wire[15:0] tmp7981;
    wire[15:0] tmp7982;
    wire[15:0] tmp7983;
    wire[15:0] tmp7984;
    wire[15:0] tmp7985;
    wire[15:0] tmp7986;
    wire[15:0] tmp7987;
    wire[15:0] tmp7988;
    wire[15:0] tmp7989;
    wire[15:0] tmp7990;
    wire[15:0] tmp7991;
    wire[15:0] tmp7992;
    wire[15:0] tmp7993;
    wire[15:0] tmp7994;
    wire[15:0] tmp7995;
    wire[15:0] tmp7996;
    wire[15:0] tmp7997;
    wire[15:0] tmp7998;
    wire[15:0] tmp7999;
    wire[15:0] tmp8000;
    wire[15:0] tmp8001;
    wire[15:0] tmp8002;
    wire tmp8003;
    wire tmp8004;
    wire tmp8005;
    wire tmp8006;
    wire tmp8007;
    wire tmp8008;
    wire tmp8009;
    wire tmp8010;
    wire tmp8011;
    wire tmp8012;
    wire tmp8013;
    wire tmp8014;
    wire tmp8015;
    wire tmp8016;
    wire tmp8017;
    wire tmp8018;
    wire[3:0] tmp8019;
    wire[3:0] tmp8020;
    wire[3:0] tmp8021;
    wire[3:0] tmp8022;
    wire[3:0] tmp8023;
    wire[3:0] tmp8024;
    wire[3:0] tmp8025;
    wire[3:0] tmp8026;
    wire[3:0] tmp8027;
    wire[3:0] tmp8028;
    wire[3:0] tmp8029;
    wire[3:0] tmp8030;
    wire[3:0] tmp8031;
    wire[3:0] tmp8032;
    wire[3:0] tmp8033;
    wire tmp8034;
    wire tmp8035;
    wire tmp8036;
    wire tmp8037;
    wire tmp8038;
    wire[15:0] tmp8041;
    wire[15:0] tmp8042;
    wire[15:0] tmp8045;
    wire[15:0] tmp8046;
    wire[15:0] tmp8049;
    wire[15:0] tmp8050;
    wire[15:0] tmp8053;
    wire[15:0] tmp8054;
    wire[15:0] tmp8057;
    wire[15:0] tmp8058;
    wire[15:0] tmp8061;
    wire[15:0] tmp8062;
    wire[15:0] tmp8065;
    wire[15:0] tmp8066;
    wire[15:0] tmp8069;
    wire[15:0] tmp8070;
    wire tmp8074;
    wire[3:0] tmp8076;
    wire tmp8077;
    wire tmp8078;
    wire[3:0] tmp8080;
    wire tmp8081;
    wire tmp8082;
    wire tmp8083;
    wire tmp8084;
    wire tmp8087;
    wire tmp8090;
    wire tmp8091;
    wire tmp8095;
    wire tmp8099;
    wire tmp8101;
    wire tmp8102;
    wire[3:0] tmp8104;
    wire tmp8105;
    wire tmp8106;
    wire[3:0] tmp8108;
    wire tmp8109;
    wire tmp8110;
    wire tmp8112;
    wire tmp8114;
    wire[2:0] tmp8117;
    wire tmp8118;
    wire tmp8120;
    wire tmp8126;
    wire tmp8129;
    wire tmp8130;
    wire tmp8138;
    wire tmp8141;
    wire tmp8144;
    wire tmp8149;
    wire tmp8156;
    wire[2:0] tmp8157;
    wire[2:0] tmp8158;
    wire[2:0] tmp8159;
    wire[2:0] tmp8160;
    wire[3:0] tmp8161;
    wire[3:0] tmp8162;
    wire[3:0] tmp8163;
    wire[3:0] tmp8164;

    // Combinational
    assign _ver_out_tmp_0 = 32768;
    assign _ver_out_tmp_1 = 32768;
    assign _ver_out_tmp_2 = 32768;
    assign _ver_out_tmp_3 = 32768;
    assign _ver_out_tmp_4 = 32768;
    assign _ver_out_tmp_5 = 32768;
    assign _ver_out_tmp_6 = 32768;
    assign _ver_out_tmp_7 = 32768;
    assign _ver_out_tmp_8 = 32768;
    assign _ver_out_tmp_9 = 32768;
    assign _ver_out_tmp_10 = 32768;
    assign _ver_out_tmp_11 = 32768;
    assign _ver_out_tmp_12 = 32768;
    assign _ver_out_tmp_13 = 32768;
    assign _ver_out_tmp_14 = 32768;
    assign _ver_out_tmp_15 = 32768;
    assign _ver_out_tmp_16 = 32768;
    assign _ver_out_tmp_17 = 32768;
    assign _ver_out_tmp_18 = 32768;
    assign _ver_out_tmp_19 = 32768;
    assign _ver_out_tmp_20 = 32768;
    assign _ver_out_tmp_21 = 32768;
    assign _ver_out_tmp_22 = 32768;
    assign _ver_out_tmp_23 = 32768;
    assign _ver_out_tmp_24 = 32768;
    assign _ver_out_tmp_25 = 32768;
    assign _ver_out_tmp_26 = 32768;
    assign _ver_out_tmp_27 = 32768;
    assign _ver_out_tmp_28 = 32768;
    assign _ver_out_tmp_29 = 32768;
    assign _ver_out_tmp_30 = 32768;
    assign _ver_out_tmp_31 = 32768;
    assign _ver_out_tmp_32 = 32768;
    assign _ver_out_tmp_33 = 32768;
    assign _ver_out_tmp_34 = 32768;
    assign _ver_out_tmp_35 = 32768;
    assign _ver_out_tmp_36 = 32768;
    assign _ver_out_tmp_37 = 32768;
    assign _ver_out_tmp_38 = 32768;
    assign _ver_out_tmp_39 = 32768;
    assign _ver_out_tmp_40 = 32768;
    assign _ver_out_tmp_41 = 32768;
    assign _ver_out_tmp_42 = 32768;
    assign _ver_out_tmp_43 = 32768;
    assign _ver_out_tmp_44 = 32768;
    assign _ver_out_tmp_45 = 32768;
    assign _ver_out_tmp_46 = 32768;
    assign _ver_out_tmp_47 = 32768;
    assign _ver_out_tmp_48 = 32768;
    assign _ver_out_tmp_49 = 32768;
    assign _ver_out_tmp_50 = 32768;
    assign _ver_out_tmp_51 = 32768;
    assign _ver_out_tmp_52 = 32768;
    assign _ver_out_tmp_53 = 32768;
    assign _ver_out_tmp_54 = 32768;
    assign _ver_out_tmp_55 = 32768;
    assign _ver_out_tmp_56 = 32768;
    assign _ver_out_tmp_57 = 32768;
    assign _ver_out_tmp_58 = 32768;
    assign _ver_out_tmp_59 = 32768;
    assign _ver_out_tmp_60 = 32768;
    assign _ver_out_tmp_61 = 32768;
    assign _ver_out_tmp_62 = 32768;
    assign _ver_out_tmp_63 = 32768;
    assign _ver_out_tmp_64 = 32768;
    assign _ver_out_tmp_65 = 32768;
    assign _ver_out_tmp_66 = 32768;
    assign _ver_out_tmp_67 = 32768;
    assign _ver_out_tmp_68 = 32768;
    assign _ver_out_tmp_69 = 32768;
    assign _ver_out_tmp_70 = 32768;
    assign _ver_out_tmp_71 = 32768;
    assign _ver_out_tmp_72 = 32768;
    assign _ver_out_tmp_73 = 32768;
    assign _ver_out_tmp_74 = 32768;
    assign _ver_out_tmp_75 = 32768;
    assign _ver_out_tmp_76 = 32768;
    assign _ver_out_tmp_77 = 32768;
    assign _ver_out_tmp_78 = 32768;
    assign _ver_out_tmp_79 = 32768;
    assign _ver_out_tmp_80 = 32768;
    assign _ver_out_tmp_81 = 32768;
    assign _ver_out_tmp_82 = 32768;
    assign _ver_out_tmp_83 = 32768;
    assign _ver_out_tmp_84 = 32768;
    assign _ver_out_tmp_85 = 32768;
    assign _ver_out_tmp_86 = 32768;
    assign _ver_out_tmp_87 = 32768;
    assign _ver_out_tmp_88 = 32768;
    assign _ver_out_tmp_89 = 32768;
    assign _ver_out_tmp_90 = 32768;
    assign _ver_out_tmp_91 = 32768;
    assign const_1_1 = 1;
    assign const_2_0 = 0;
    assign const_3_0 = 0;
    assign const_4_0 = 0;
    assign const_5_4 = 4;
    assign const_6_0 = 0;
    assign const_7_2 = 2;
    assign const_8_1 = 1;
    assign const_9_0 = 0;
    assign const_10_0 = 0;
    assign const_11_0 = 0;
    assign const_12_0 = 0;
    assign const_13_1 = 1;
    assign const_14_0 = 0;
    assign const_15_1 = 1;
    assign const_16_0 = 0;
    assign const_17_0 = 0;
    assign const_18_0 = 0;
    assign const_19_0 = 0;
    assign const_20_15 = 15;
    assign const_21_1 = 1;
    assign const_22_0 = 0;
    assign const_23_2 = 2;
    assign const_24_0 = 0;
    assign const_25_3 = 3;
    assign const_26_0 = 0;
    assign const_27_0 = 0;
    assign const_28_0 = 0;
    assign const_29_0 = 0;
    assign const_30_0 = 0;
    assign const_31_0 = 0;
    assign const_32_32767 = 32767;
    assign const_34_0 = 0;
    assign const_35_0 = 0;
    assign const_36_0 = 0;
    assign const_37_0 = 0;
    assign const_38_0 = 0;
    assign const_39_32767 = 32767;
    assign const_41_0 = 0;
    assign const_42_0 = 0;
    assign const_43_0 = 0;
    assign const_44_0 = 0;
    assign const_45_0 = 0;
    assign const_46_32767 = 32767;
    assign const_48_0 = 0;
    assign const_49_0 = 0;
    assign const_50_0 = 0;
    assign const_51_0 = 0;
    assign const_52_0 = 0;
    assign const_53_32767 = 32767;
    assign const_55_6 = 6;
    assign const_56_0 = 0;
    assign const_57_7 = 7;
    assign const_58_0 = 0;
    assign const_59_4 = 4;
    assign const_60_0 = 0;
    assign const_61_5 = 5;
    assign const_62_0 = 0;
    assign const_63_0 = 0;
    assign const_64_0 = 0;
    assign const_65_0 = 0;
    assign const_66_0 = 0;
    assign const_67_0 = 0;
    assign const_68_0 = 0;
    assign const_69_32767 = 32767;
    assign const_71_0 = 0;
    assign const_72_0 = 0;
    assign const_73_0 = 0;
    assign const_74_0 = 0;
    assign const_75_0 = 0;
    assign const_76_0 = 0;
    assign const_77_32767 = 32767;
    assign const_79_0 = 0;
    assign const_80_0 = 0;
    assign const_81_0 = 0;
    assign const_82_0 = 0;
    assign const_83_0 = 0;
    assign const_84_0 = 0;
    assign const_85_32767 = 32767;
    assign const_87_0 = 0;
    assign const_88_0 = 0;
    assign const_89_0 = 0;
    assign const_90_0 = 0;
    assign const_91_0 = 0;
    assign const_92_0 = 0;
    assign const_93_32767 = 32767;
    assign const_95_8 = 8;
    assign const_97_0 = 0;
    assign const_98_0 = 0;
    assign const_99_32767 = 32767;
    assign const_100_0 = 0;
    assign const_102_0 = 0;
    assign const_103_0 = 0;
    assign const_104_32767 = 32767;
    assign const_105_0 = 0;
    assign const_107_0 = 0;
    assign const_108_0 = 0;
    assign const_109_32767 = 32767;
    assign const_110_0 = 0;
    assign const_112_0 = 0;
    assign const_113_0 = 0;
    assign const_114_32767 = 32767;
    assign const_115_0 = 0;
    assign const_116_2 = 2;
    assign const_117_0 = 0;
    assign const_118_0 = 0;
    assign const_119_0 = 0;
    assign const_120_0 = 0;
    assign const_121_15 = 15;
    assign const_122_1 = 1;
    assign const_123_0 = 0;
    assign const_124_2 = 2;
    assign const_125_0 = 0;
    assign const_126_3 = 3;
    assign const_127_0 = 0;
    assign const_128_0 = 0;
    assign const_129_0 = 0;
    assign const_130_0 = 0;
    assign const_131_0 = 0;
    assign const_132_0 = 0;
    assign const_133_32767 = 32767;
    assign const_135_0 = 0;
    assign const_136_0 = 0;
    assign const_137_0 = 0;
    assign const_138_0 = 0;
    assign const_139_0 = 0;
    assign const_140_32767 = 32767;
    assign const_142_0 = 0;
    assign const_143_0 = 0;
    assign const_144_0 = 0;
    assign const_145_0 = 0;
    assign const_146_0 = 0;
    assign const_147_32767 = 32767;
    assign const_149_0 = 0;
    assign const_150_0 = 0;
    assign const_151_0 = 0;
    assign const_152_0 = 0;
    assign const_153_0 = 0;
    assign const_154_32767 = 32767;
    assign const_156_6 = 6;
    assign const_157_0 = 0;
    assign const_158_7 = 7;
    assign const_159_0 = 0;
    assign const_160_4 = 4;
    assign const_161_0 = 0;
    assign const_162_5 = 5;
    assign const_163_0 = 0;
    assign const_164_0 = 0;
    assign const_165_0 = 0;
    assign const_166_0 = 0;
    assign const_167_0 = 0;
    assign const_168_0 = 0;
    assign const_169_0 = 0;
    assign const_170_32767 = 32767;
    assign const_172_0 = 0;
    assign const_173_0 = 0;
    assign const_174_0 = 0;
    assign const_175_0 = 0;
    assign const_176_0 = 0;
    assign const_177_0 = 0;
    assign const_178_32767 = 32767;
    assign const_180_0 = 0;
    assign const_181_0 = 0;
    assign const_182_0 = 0;
    assign const_183_0 = 0;
    assign const_184_0 = 0;
    assign const_185_0 = 0;
    assign const_186_32767 = 32767;
    assign const_188_0 = 0;
    assign const_189_0 = 0;
    assign const_190_0 = 0;
    assign const_191_0 = 0;
    assign const_192_0 = 0;
    assign const_193_0 = 0;
    assign const_194_32767 = 32767;
    assign const_196_8 = 8;
    assign const_198_0 = 0;
    assign const_199_0 = 0;
    assign const_200_32767 = 32767;
    assign const_201_0 = 0;
    assign const_203_0 = 0;
    assign const_204_0 = 0;
    assign const_205_32767 = 32767;
    assign const_206_0 = 0;
    assign const_208_0 = 0;
    assign const_209_0 = 0;
    assign const_210_32767 = 32767;
    assign const_211_0 = 0;
    assign const_213_0 = 0;
    assign const_214_0 = 0;
    assign const_215_32767 = 32767;
    assign const_216_0 = 0;
    assign const_217_3 = 3;
    assign const_218_0 = 0;
    assign const_219_0 = 0;
    assign const_220_0 = 0;
    assign const_221_0 = 0;
    assign const_222_0 = 0;
    assign const_223_0 = 0;
    assign const_224_0 = 0;
    assign const_225_0 = 0;
    assign const_226_0 = 0;
    assign const_227_0 = 0;
    assign const_228_0 = 0;
    assign const_229_0 = 0;
    assign const_230_0 = 0;
    assign const_231_0 = 0;
    assign const_232_0 = 0;
    assign const_233_0 = 0;
    assign const_234_0 = 0;
    assign const_235_0 = 0;
    assign const_236_0 = 0;
    assign const_237_0 = 0;
    assign const_238_0 = 0;
    assign const_239_0 = 0;
    assign const_240_0 = 0;
    assign const_242_0 = 0;
    assign const_243_0 = 0;
    assign const_244_32767 = 32767;
    assign const_245_0 = 0;
    assign const_247_0 = 0;
    assign const_248_0 = 0;
    assign const_249_32767 = 32767;
    assign const_250_0 = 0;
    assign const_252_0 = 0;
    assign const_253_0 = 0;
    assign const_254_32767 = 32767;
    assign const_255_0 = 0;
    assign const_257_0 = 0;
    assign const_258_0 = 0;
    assign const_259_32767 = 32767;
    assign const_260_0 = 0;
    assign const_262_0 = 0;
    assign const_263_0 = 0;
    assign const_264_32767 = 32767;
    assign const_265_0 = 0;
    assign const_267_0 = 0;
    assign const_268_0 = 0;
    assign const_269_32767 = 32767;
    assign const_270_0 = 0;
    assign const_272_0 = 0;
    assign const_273_0 = 0;
    assign const_274_32767 = 32767;
    assign const_275_0 = 0;
    assign const_277_0 = 0;
    assign const_278_0 = 0;
    assign const_279_32767 = 32767;
    assign const_280_0 = 0;
    assign const_281_0 = 0;
    assign const_282_0 = 0;
    assign const_283_0 = 0;
    assign const_284_0 = 0;
    assign const_285_0 = 0;
    assign const_286_0 = 0;
    assign const_287_0 = 0;
    assign const_288_0 = 0;
    assign const_289_0 = 0;
    assign const_290_0 = 0;
    assign const_291_15 = 15;
    assign const_292_0 = 0;
    assign const_293_0 = 0;
    assign const_294_0 = 0;
    assign const_295_8 = 8;
    assign const_296_0 = 0;
    assign const_298_0 = 0;
    assign const_299_0 = 0;
    assign const_300_32767 = 32767;
    assign const_301_0 = 0;
    assign const_303_0 = 0;
    assign const_304_0 = 0;
    assign const_305_32767 = 32767;
    assign const_306_0 = 0;
    assign const_308_0 = 0;
    assign const_309_0 = 0;
    assign const_310_32767 = 32767;
    assign const_311_0 = 0;
    assign const_313_0 = 0;
    assign const_314_0 = 0;
    assign const_315_32767 = 32767;
    assign const_316_0 = 0;
    assign const_317_1 = 1;
    assign const_318_0 = 0;
    assign const_319_0 = 0;
    assign const_320_0 = 0;
    assign const_321_0 = 0;
    assign const_322_0 = 0;
    assign const_323_0 = 0;
    assign const_324_32767 = 32767;
    assign const_326_0 = 0;
    assign const_327_0 = 0;
    assign const_328_0 = 0;
    assign const_329_0 = 0;
    assign const_330_0 = 0;
    assign const_331_32767 = 32767;
    assign const_333_0 = 0;
    assign const_334_0 = 0;
    assign const_335_0 = 0;
    assign const_336_0 = 0;
    assign const_337_0 = 0;
    assign const_338_32767 = 32767;
    assign const_340_0 = 0;
    assign const_341_0 = 0;
    assign const_342_0 = 0;
    assign const_343_0 = 0;
    assign const_344_0 = 0;
    assign const_345_32767 = 32767;
    assign const_347_4 = 4;
    assign const_348_0 = 0;
    assign const_350_0 = 0;
    assign const_351_0 = 0;
    assign const_352_32767 = 32767;
    assign const_353_0 = 0;
    assign const_354_0 = 0;
    assign const_355_0 = 0;
    assign const_356_0 = 0;
    assign const_357_0 = 0;
    assign const_358_0 = 0;
    assign const_359_0 = 0;
    assign const_360_32767 = 32767;
    assign const_363_0 = 0;
    assign const_364_0 = 0;
    assign const_365_32767 = 32767;
    assign const_366_0 = 0;
    assign const_367_0 = 0;
    assign const_368_0 = 0;
    assign const_369_0 = 0;
    assign const_370_0 = 0;
    assign const_371_0 = 0;
    assign const_372_0 = 0;
    assign const_373_32767 = 32767;
    assign const_376_0 = 0;
    assign const_377_0 = 0;
    assign const_378_32767 = 32767;
    assign const_379_0 = 0;
    assign const_380_0 = 0;
    assign const_381_0 = 0;
    assign const_382_0 = 0;
    assign const_383_0 = 0;
    assign const_384_0 = 0;
    assign const_385_0 = 0;
    assign const_386_32767 = 32767;
    assign const_389_0 = 0;
    assign const_390_0 = 0;
    assign const_391_32767 = 32767;
    assign const_392_0 = 0;
    assign const_393_0 = 0;
    assign const_394_0 = 0;
    assign const_395_0 = 0;
    assign const_396_0 = 0;
    assign const_397_0 = 0;
    assign const_398_0 = 0;
    assign const_399_32767 = 32767;
    assign const_401_6 = 6;
    assign const_402_0 = 0;
    assign const_403_0 = 0;
    assign const_404_0 = 0;
    assign const_405_0 = 0;
    assign const_406_0 = 0;
    assign const_407_0 = 0;
    assign const_408_32767 = 32767;
    assign const_410_0 = 0;
    assign const_411_0 = 0;
    assign const_412_0 = 0;
    assign const_413_0 = 0;
    assign const_414_0 = 0;
    assign const_415_32767 = 32767;
    assign const_417_0 = 0;
    assign const_418_0 = 0;
    assign const_419_0 = 0;
    assign const_420_0 = 0;
    assign const_421_0 = 0;
    assign const_422_32767 = 32767;
    assign const_424_0 = 0;
    assign const_425_0 = 0;
    assign const_426_0 = 0;
    assign const_427_0 = 0;
    assign const_428_0 = 0;
    assign const_429_32767 = 32767;
    assign const_431_2 = 2;
    assign const_432_0 = 0;
    assign const_433_0 = 0;
    assign const_434_0 = 0;
    assign const_435_0 = 0;
    assign const_436_0 = 0;
    assign const_437_0 = 0;
    assign const_438_32767 = 32767;
    assign const_440_0 = 0;
    assign const_441_0 = 0;
    assign const_442_0 = 0;
    assign const_443_0 = 0;
    assign const_444_0 = 0;
    assign const_445_32767 = 32767;
    assign const_447_0 = 0;
    assign const_448_0 = 0;
    assign const_449_0 = 0;
    assign const_450_0 = 0;
    assign const_451_0 = 0;
    assign const_452_32767 = 32767;
    assign const_454_0 = 0;
    assign const_455_0 = 0;
    assign const_456_0 = 0;
    assign const_457_0 = 0;
    assign const_458_0 = 0;
    assign const_459_32767 = 32767;
    assign const_461_0 = 0;
    assign const_462_0 = 0;
    assign const_463_0 = 0;
    assign const_464_0 = 0;
    assign const_465_0 = 0;
    assign const_466_32767 = 32767;
    assign const_468_0 = 0;
    assign const_469_0 = 0;
    assign const_470_0 = 0;
    assign const_471_0 = 0;
    assign const_472_0 = 0;
    assign const_473_32767 = 32767;
    assign const_475_0 = 0;
    assign const_476_0 = 0;
    assign const_477_0 = 0;
    assign const_478_0 = 0;
    assign const_479_0 = 0;
    assign const_480_32767 = 32767;
    assign const_482_0 = 0;
    assign const_483_0 = 0;
    assign const_484_0 = 0;
    assign const_485_0 = 0;
    assign const_486_0 = 0;
    assign const_487_32767 = 32767;
    assign const_489_0 = 0;
    assign const_490_0 = 0;
    assign const_491_0 = 0;
    assign const_492_0 = 0;
    assign const_493_0 = 0;
    assign const_494_32767 = 32767;
    assign const_496_0 = 0;
    assign const_497_0 = 0;
    assign const_498_0 = 0;
    assign const_499_0 = 0;
    assign const_500_0 = 0;
    assign const_501_32767 = 32767;
    assign const_503_0 = 0;
    assign const_504_0 = 0;
    assign const_505_0 = 0;
    assign const_506_0 = 0;
    assign const_507_0 = 0;
    assign const_508_32767 = 32767;
    assign const_510_0 = 0;
    assign const_511_0 = 0;
    assign const_512_0 = 0;
    assign const_513_0 = 0;
    assign const_514_0 = 0;
    assign const_515_32767 = 32767;
    assign const_517_5 = 5;
    assign const_518_1 = 1;
    assign const_520_0 = 0;
    assign const_521_0 = 0;
    assign const_522_32767 = 32767;
    assign const_523_0 = 0;
    assign const_524_0 = 0;
    assign const_525_0 = 0;
    assign const_526_0 = 0;
    assign const_527_0 = 0;
    assign const_528_0 = 0;
    assign const_529_0 = 0;
    assign const_530_32767 = 32767;
    assign const_533_0 = 0;
    assign const_534_0 = 0;
    assign const_535_32767 = 32767;
    assign const_536_0 = 0;
    assign const_537_0 = 0;
    assign const_538_0 = 0;
    assign const_539_0 = 0;
    assign const_540_0 = 0;
    assign const_541_0 = 0;
    assign const_542_0 = 0;
    assign const_543_32767 = 32767;
    assign const_546_0 = 0;
    assign const_547_0 = 0;
    assign const_548_32767 = 32767;
    assign const_549_0 = 0;
    assign const_550_0 = 0;
    assign const_551_0 = 0;
    assign const_552_0 = 0;
    assign const_553_0 = 0;
    assign const_554_0 = 0;
    assign const_555_0 = 0;
    assign const_556_32767 = 32767;
    assign const_559_0 = 0;
    assign const_560_0 = 0;
    assign const_561_32767 = 32767;
    assign const_562_0 = 0;
    assign const_563_0 = 0;
    assign const_564_0 = 0;
    assign const_565_0 = 0;
    assign const_566_0 = 0;
    assign const_567_0 = 0;
    assign const_568_0 = 0;
    assign const_569_32767 = 32767;
    assign const_571_0 = 0;
    assign const_572_0 = 0;
    assign const_573_0 = 0;
    assign const_574_0 = 0;
    assign const_575_0 = 0;
    assign const_577_0 = 0;
    assign const_578_0 = 0;
    assign const_579_32767 = 32767;
    assign const_580_0 = 0;
    assign const_581_0 = 0;
    assign const_582_0 = 0;
    assign const_584_0 = 0;
    assign const_585_0 = 0;
    assign const_586_32767 = 32767;
    assign const_587_0 = 0;
    assign const_588_0 = 0;
    assign const_589_0 = 0;
    assign const_591_0 = 0;
    assign const_592_0 = 0;
    assign const_593_32767 = 32767;
    assign const_594_0 = 0;
    assign const_595_0 = 0;
    assign const_596_0 = 0;
    assign const_598_0 = 0;
    assign const_599_0 = 0;
    assign const_600_32767 = 32767;
    assign const_601_0 = 0;
    assign const_602_0 = 0;
    assign const_603_0 = 0;
    assign const_605_0 = 0;
    assign const_606_0 = 0;
    assign const_607_32767 = 32767;
    assign const_608_0 = 0;
    assign const_609_0 = 0;
    assign const_610_0 = 0;
    assign const_612_0 = 0;
    assign const_613_0 = 0;
    assign const_614_32767 = 32767;
    assign const_615_0 = 0;
    assign const_616_0 = 0;
    assign const_617_0 = 0;
    assign const_619_0 = 0;
    assign const_620_0 = 0;
    assign const_621_32767 = 32767;
    assign const_622_0 = 0;
    assign const_623_0 = 0;
    assign const_624_0 = 0;
    assign const_626_0 = 0;
    assign const_627_0 = 0;
    assign const_628_32767 = 32767;
    assign const_629_0 = 0;
    assign const_630_0 = 0;
    assign const_631_6 = 6;
    assign const_632_1 = 1;
    assign const_633_0 = 0;
    assign const_635_0 = 0;
    assign const_636_0 = 0;
    assign const_637_32767 = 32767;
    assign const_638_0 = 0;
    assign const_639_0 = 0;
    assign const_640_0 = 0;
    assign const_642_0 = 0;
    assign const_643_0 = 0;
    assign const_644_32767 = 32767;
    assign const_645_0 = 0;
    assign const_646_0 = 0;
    assign const_647_0 = 0;
    assign const_649_0 = 0;
    assign const_650_0 = 0;
    assign const_651_32767 = 32767;
    assign const_652_0 = 0;
    assign const_653_0 = 0;
    assign const_654_0 = 0;
    assign const_656_0 = 0;
    assign const_657_0 = 0;
    assign const_658_32767 = 32767;
    assign const_659_0 = 0;
    assign const_660_0 = 0;
    assign const_661_0 = 0;
    assign const_663_0 = 0;
    assign const_664_0 = 0;
    assign const_665_32767 = 32767;
    assign const_666_0 = 0;
    assign const_667_0 = 0;
    assign const_668_0 = 0;
    assign const_670_0 = 0;
    assign const_671_0 = 0;
    assign const_672_32767 = 32767;
    assign const_673_0 = 0;
    assign const_674_0 = 0;
    assign const_675_0 = 0;
    assign const_677_0 = 0;
    assign const_678_0 = 0;
    assign const_679_32767 = 32767;
    assign const_680_0 = 0;
    assign const_681_0 = 0;
    assign const_682_0 = 0;
    assign const_684_0 = 0;
    assign const_685_0 = 0;
    assign const_686_32767 = 32767;
    assign const_687_0 = 0;
    assign const_688_0 = 0;
    assign const_689_3 = 3;
    assign const_690_1 = 1;
    assign const_691_0 = 0;
    assign const_692_0 = 0;
    assign const_693_0 = 0;
    assign const_694_0 = 0;
    assign const_695_0 = 0;
    assign const_696_32767 = 32767;
    assign const_698_0 = 0;
    assign const_699_0 = 0;
    assign const_700_0 = 0;
    assign const_701_0 = 0;
    assign const_702_0 = 0;
    assign const_703_32767 = 32767;
    assign const_705_0 = 0;
    assign const_706_0 = 0;
    assign const_707_0 = 0;
    assign const_708_0 = 0;
    assign const_709_0 = 0;
    assign const_710_32767 = 32767;
    assign const_712_0 = 0;
    assign const_713_0 = 0;
    assign const_714_0 = 0;
    assign const_715_0 = 0;
    assign const_716_0 = 0;
    assign const_717_32767 = 32767;
    assign const_719_0 = 0;
    assign const_720_0 = 0;
    assign const_721_0 = 0;
    assign const_722_0 = 0;
    assign const_723_0 = 0;
    assign const_724_0 = 0;
    assign const_725_0 = 0;
    assign const_726_0 = 0;
    assign const_727_0 = 0;
    assign const_728_0 = 0;
    assign const_729_0 = 0;
    assign const_730_0 = 0;
    assign const_731_0 = 0;
    assign const_732_0 = 0;
    assign const_733_0 = 0;
    assign const_734_0 = 0;
    assign const_735_0 = 0;
    assign const_736_0 = 0;
    assign const_737_0 = 0;
    assign const_738_0 = 0;
    assign const_739_0 = 0;
    assign const_740_0 = 0;
    assign const_741_0 = 0;
    assign const_742_1 = 1;
    assign const_743_0 = 0;
    assign const_744_2 = 2;
    assign const_745_0 = 0;
    assign const_746_3 = 3;
    assign const_747_0 = 0;
    assign const_748_15 = 15;
    assign const_749_4 = 4;
    assign const_750_0 = 0;
    assign const_751_5 = 5;
    assign const_752_0 = 0;
    assign const_753_6 = 6;
    assign const_754_0 = 0;
    assign const_755_7 = 7;
    assign const_756_0 = 0;
    assign const_757_15 = 15;
    assign const_758_8 = 8;
    assign const_759_6 = 6;
    assign const_760_0 = 0;
    assign const_761_7 = 7;
    assign const_762_0 = 0;
    assign const_763_15 = 15;
    assign const_764_1 = 1;
    assign const_765_0 = 0;
    assign const_766_2 = 2;
    assign const_767_15 = 15;
    assign const_768_2 = 2;
    assign const_769_0 = 0;
    assign const_770_3 = 3;
    assign const_771_3 = 3;
    assign const_772_0 = 0;
    assign const_773_1 = 1;
    assign const_774_15 = 15;
    assign const_775_1 = 1;
    assign const_776_15 = 15;
    assign const_781_0 = 0;
    assign const_782_0 = 0;
    assign const_783_0 = 0;
    assign const_784_0 = 0;
    assign blue_o = tmp8112;
    assign green_o = tmp8101;
    assign red_o = tmp8084;
    assign tmp1 = {const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0, const_2_0};
    assign tmp2 = {tmp1, const_1_1};
    assign tmp3 = tmp0 + tmp2;
    assign tmp4 = {tmp3[26], tmp3[25], tmp3[24], tmp3[23], tmp3[22], tmp3[21], tmp3[20], tmp3[19], tmp3[18], tmp3[17], tmp3[16], tmp3[15], tmp3[14], tmp3[13], tmp3[12], tmp3[11], tmp3[10], tmp3[9], tmp3[8], tmp3[7], tmp3[6], tmp3[5], tmp3[4], tmp3[3], tmp3[2], tmp3[1], tmp3[0]};
    assign tmp8 = {tmp0[26]};
    assign tmp10 = ~tmp8114;
    assign tmp33 = ~tmp7;
    assign tmp35 = {tmp6808, const_3_0};
    assign tmp36 = my_calculator_ctrl == tmp35;
    assign tmp37 = my_calculator_ctrl == const_5_4;
    assign tmp73 = tmp2610 & tmp37;
    assign tmp90 = {tmp1178, const_18_0};
    assign tmp91 = my_calculator_in_x == tmp90;
    assign tmp92 = my_calculator_in_x == const_20_15;
    assign tmp119 = tmp1051 & tmp92;
    assign tmp131 = my_calculator_in_x == tmp1179;
    assign tmp134 = my_calculator_in_x == tmp8076;
    assign tmp135 = tmp131 | tmp134;
    assign tmp138 = my_calculator_in_x == tmp8080;
    assign tmp139 = tmp135 | tmp138;
    assign tmp141 = {tmp1189, const_27_0};
    assign tmp143 = {const_28_0, const_28_0, const_28_0, const_28_0, const_28_0, const_28_0, const_28_0, const_28_0, const_28_0, const_28_0, const_28_0, const_28_0, const_28_0, const_28_0, const_28_0};
    assign tmp150 = tmp1196 ^ tmp6605;
    assign tmp152 = ~tmp2625;
    assign tmp158 = tmp141 - tmp2887;
    assign tmp160 = {tmp141[15]};
    assign tmp161 = ~tmp160;
    assign tmp162 = tmp1208 ^ tmp161;
    assign tmp166 = tmp1202 & tmp1214;
    assign tmp183 = tmp2887 - tmp141;
    assign tmp190 = tmp1236 ^ tmp161;
    assign tmp192 = tmp190 | tmp1240;
    assign tmp193 = tmp586 & tmp192;
    assign tmp194 = tmp166 ? const_32_32767 : tmp141;
    assign tmp195 = tmp193 ? _ver_out_tmp_14 : tmp194;
    assign tmp207 = {tmp12[14], tmp12[13], tmp12[12], tmp12[11], tmp12[10], tmp12[9], tmp12[8], tmp12[7], tmp12[6], tmp12[5], tmp12[4], tmp12[3], tmp12[2], tmp12[1], tmp12[0]};
    assign tmp208 = {tmp207, const_34_0};
    assign tmp217 = tmp1625 ^ tmp6605;
    assign tmp225 = tmp208 - tmp2887;
    assign tmp226 = {tmp225[16]};
    assign tmp228 = ~tmp255;
    assign tmp229 = tmp226 ^ tmp228;
    assign tmp232 = tmp229 ^ tmp6605;
    assign tmp233 = tmp667 & tmp232;
    assign tmp250 = tmp2887 - tmp208;
    assign tmp251 = {tmp250[16]};
    assign tmp254 = tmp251 ^ tmp6605;
    assign tmp255 = {tmp208[15]};
    assign tmp257 = tmp254 ^ tmp228;
    assign tmp258 = tmp2887 == tmp208;
    assign tmp259 = tmp257 | tmp258;
    assign tmp260 = tmp2247 & tmp259;
    assign tmp261 = tmp233 ? const_39_32767 : tmp208;
    assign tmp262 = tmp260 ? _ver_out_tmp_17 : tmp261;
    assign tmp269 = ~tmp91;
    assign tmp273 = tmp424 & tmp139;
    assign tmp274 = {tmp15[14], tmp15[13], tmp15[12], tmp15[11], tmp15[10], tmp15[9], tmp15[8], tmp15[7], tmp15[6], tmp15[5], tmp15[4], tmp15[3], tmp15[2], tmp15[1], tmp15[0]};
    assign tmp292 = tmp1328 - tmp2887;
    assign tmp293 = {tmp292[16]};
    assign tmp318 = {tmp1370[16]};
    assign tmp321 = tmp318 ^ tmp6605;
    assign tmp325 = tmp2887 == tmp1328;
    assign tmp329 = tmp1380 ? _ver_out_tmp_21 : tmp1381;
    assign tmp342 = {tmp7565, const_48_0};
    assign tmp351 = tmp7572 ^ tmp6605;
    assign tmp354 = tmp351 ^ tmp7577;
    assign tmp359 = tmp342 - tmp2887;
    assign tmp360 = {tmp359[16]};
    assign tmp362 = ~tmp389;
    assign tmp376 = tmp943 ^ tmp7577;
    assign tmp384 = tmp2887 - tmp342;
    assign tmp385 = {tmp384[16]};
    assign tmp388 = tmp385 ^ tmp6605;
    assign tmp389 = {tmp342[15]};
    assign tmp392 = tmp2887 == tmp342;
    assign tmp395 = tmp7591 ? const_53_32767 : tmp342;
    assign tmp410 = my_calculator_in_x == tmp8104;
    assign tmp413 = my_calculator_in_x == tmp8108;
    assign tmp414 = tmp410 | tmp413;
    assign tmp423 = ~tmp92;
    assign tmp424 = tmp1051 & tmp423;
    assign tmp427 = tmp764 & tmp414;
    assign tmp459 = tmp4971 & tmp8118;
    assign tmp520 = {const_60_0, const_59_4};
    assign tmp521 = my_calculator_in_x == tmp520;
    assign tmp523 = {const_62_0, const_61_5};
    assign tmp524 = my_calculator_in_x == tmp523;
    assign tmp525 = tmp521 | tmp524;
    assign tmp532 = tmp1601 + tmp1726;
    assign tmp533 = {tmp532[16], tmp532[15], tmp532[14], tmp532[13], tmp532[12], tmp532[11], tmp532[10], tmp532[9], tmp532[8], tmp532[7], tmp532[6], tmp532[5], tmp532[4], tmp532[3], tmp532[2], tmp532[1], tmp532[0]};
    assign tmp534 = {tmp533[15], tmp533[14], tmp533[13], tmp533[12], tmp533[11], tmp533[10], tmp533[9], tmp533[8], tmp533[7], tmp533[6], tmp533[5], tmp533[4], tmp533[3], tmp533[2], tmp533[1], tmp533[0]};
    assign tmp558 = tmp1268 ^ tmp1743;
    assign tmp559 = tmp1202 & tmp558;
    assign tmp564 = tmp534 - tmp2887;
    assign tmp565 = {tmp564[16]};
    assign tmp566 = {tmp534[15]};
    assign tmp568 = tmp565 ^ tmp610;
    assign tmp571 = tmp568 ^ tmp6605;
    assign tmp573 = tmp571 | tmp612;
    assign tmp574 = tmp559 & tmp573;
    assign tmp579 = tmp11 - tmp2887;
    assign tmp586 = tmp2627 ^ tmp6605;
    assign tmp592 = {tmp6851[16]};
    assign tmp593 = {tmp13[15]};
    assign tmp595 = tmp592 ^ tmp1743;
    assign tmp599 = tmp586 & tmp7250;
    assign tmp604 = tmp2887 - tmp534;
    assign tmp605 = {tmp604[16]};
    assign tmp608 = tmp605 ^ tmp6605;
    assign tmp610 = ~tmp566;
    assign tmp611 = tmp608 ^ tmp610;
    assign tmp612 = tmp2887 == tmp534;
    assign tmp613 = tmp611 | tmp612;
    assign tmp614 = tmp599 & tmp613;
    assign tmp615 = tmp574 ? const_69_32767 : tmp534;
    assign tmp616 = tmp614 ? _ver_out_tmp_30 : tmp615;
    assign tmp642 = ~tmp139;
    assign tmp650 = {tmp14[15]};
    assign tmp653 = tmp1604 + tmp1729;
    assign tmp654 = {tmp653[16], tmp653[15], tmp653[14], tmp653[13], tmp653[12], tmp653[11], tmp653[10], tmp653[9], tmp653[8], tmp653[7], tmp653[6], tmp653[5], tmp653[4], tmp653[3], tmp653[2], tmp653[1], tmp653[0]};
    assign tmp655 = {tmp654[15], tmp654[14], tmp654[13], tmp654[12], tmp654[11], tmp654[10], tmp654[9], tmp654[8], tmp654[7], tmp654[6], tmp654[5], tmp654[4], tmp654[3], tmp654[2], tmp654[1], tmp654[0]};
    assign tmp667 = tmp217 ^ tmp7185;
    assign tmp679 = tmp1753 ^ tmp2281;
    assign tmp680 = tmp667 & tmp679;
    assign tmp685 = tmp655 - tmp2887;
    assign tmp686 = {tmp685[16]};
    assign tmp689 = tmp686 ^ tmp731;
    assign tmp692 = tmp689 ^ tmp6605;
    assign tmp693 = tmp655 == tmp2887;
    assign tmp694 = tmp692 | tmp693;
    assign tmp695 = tmp680 & tmp694;
    assign tmp720 = tmp2247 & tmp6913;
    assign tmp725 = tmp2887 - tmp655;
    assign tmp726 = {tmp725[16]};
    assign tmp729 = tmp726 ^ tmp6605;
    assign tmp730 = {tmp655[15]};
    assign tmp731 = ~tmp730;
    assign tmp732 = tmp729 ^ tmp731;
    assign tmp734 = tmp732 | tmp693;
    assign tmp735 = tmp720 & tmp734;
    assign tmp736 = tmp695 ? const_77_32767 : tmp655;
    assign tmp737 = tmp735 ? _ver_out_tmp_34 : tmp736;
    assign tmp764 = tmp424 & tmp642;
    assign tmp770 = {tmp1849, tmp15};
    assign tmp774 = tmp770 + tmp1976;
    assign tmp775 = {tmp774[16], tmp774[15], tmp774[14], tmp774[13], tmp774[12], tmp774[11], tmp774[10], tmp774[9], tmp774[8], tmp774[7], tmp774[6], tmp774[5], tmp774[4], tmp774[3], tmp774[2], tmp774[1], tmp774[0]};
    assign tmp776 = {tmp775[15], tmp775[14], tmp775[13], tmp775[12], tmp775[11], tmp775[10], tmp775[9], tmp775[8], tmp775[7], tmp775[6], tmp775[5], tmp775[4], tmp775[3], tmp775[2], tmp775[1], tmp775[0]};
    assign tmp782 = {tmp7495[16]};
    assign tmp801 = tmp1340 & tmp7654;
    assign tmp806 = tmp776 - tmp2887;
    assign tmp807 = {tmp806[16]};
    assign tmp810 = tmp807 ^ tmp852;
    assign tmp813 = tmp810 ^ tmp6605;
    assign tmp814 = tmp776 == tmp2887;
    assign tmp815 = tmp813 | tmp814;
    assign tmp816 = tmp801 & tmp815;
    assign tmp834 = {tmp2353[16]};
    assign tmp841 = tmp7154 & tmp2034;
    assign tmp846 = tmp2887 - tmp776;
    assign tmp847 = {tmp846[16]};
    assign tmp850 = tmp847 ^ tmp6605;
    assign tmp851 = {tmp776[15]};
    assign tmp852 = ~tmp851;
    assign tmp853 = tmp850 ^ tmp852;
    assign tmp855 = tmp853 | tmp814;
    assign tmp856 = tmp841 & tmp855;
    assign tmp857 = tmp816 ? const_85_32767 : tmp776;
    assign tmp858 = tmp856 ? _ver_out_tmp_37 : tmp857;
    assign tmp873 = tmp1057 & tmp525;
    assign tmp889 = {tmp16[15]};
    assign tmp895 = tmp1854 + tmp1979;
    assign tmp896 = {tmp895[16], tmp895[15], tmp895[14], tmp895[13], tmp895[12], tmp895[11], tmp895[10], tmp895[9], tmp895[8], tmp895[7], tmp895[6], tmp895[5], tmp895[4], tmp895[3], tmp895[2], tmp895[1], tmp895[0]};
    assign tmp897 = {tmp896[15], tmp896[14], tmp896[13], tmp896[12], tmp896[11], tmp896[10], tmp896[9], tmp896[8], tmp896[7], tmp896[6], tmp896[5], tmp896[4], tmp896[3], tmp896[2], tmp896[1], tmp896[0]};
    assign tmp915 = {tmp1999[16]};
    assign tmp918 = tmp915 ^ tmp6605;
    assign tmp922 = tmp354 & tmp2006;
    assign tmp927 = tmp897 - tmp2887;
    assign tmp928 = {tmp927[16]};
    assign tmp929 = {tmp897[15]};
    assign tmp930 = ~tmp929;
    assign tmp931 = tmp928 ^ tmp930;
    assign tmp934 = tmp931 ^ tmp6605;
    assign tmp935 = tmp897 == tmp2887;
    assign tmp936 = tmp934 | tmp935;
    assign tmp937 = tmp922 & tmp936;
    assign tmp943 = {tmp7596[16]};
    assign tmp962 = tmp6825 & tmp6935;
    assign tmp967 = tmp2887 - tmp897;
    assign tmp968 = {tmp967[16]};
    assign tmp971 = tmp968 ^ tmp6605;
    assign tmp974 = tmp971 ^ tmp930;
    assign tmp976 = tmp974 | tmp935;
    assign tmp977 = tmp962 & tmp976;
    assign tmp978 = tmp937 ? const_93_32767 : tmp897;
    assign tmp979 = tmp977 ? _ver_out_tmp_76 : tmp978;
    assign tmp1010 = my_calculator_in_x == const_95_8;
    assign tmp1051 = tmp459 & tmp269;
    assign tmp1057 = tmp764 & tmp1106;
    assign tmp1083 = ~tmp525;
    assign tmp1086 = tmp16 == _ver_out_tmp_47;
    assign tmp1092 = tmp1086 ? tmp6864 : tmp2565;
    assign tmp1106 = ~tmp414;
    assign tmp1109 = tmp1057 & tmp1083;
    assign tmp1110 = tmp1109 & tmp1010;
    assign tmp1112 = {const_117_0, const_116_2};
    assign tmp1113 = my_calculator_ctrl == tmp1112;
    assign tmp1132 = my_calculator_in_y == tmp90;
    assign tmp1133 = my_calculator_in_y == const_121_15;
    assign tmp1141 = tmp7818 & tmp1113;
    assign tmp1166 = tmp1841 & tmp1133;
    assign tmp1178 = {const_123_0, const_123_0, const_123_0};
    assign tmp1179 = {tmp1178, const_122_1};
    assign tmp1180 = my_calculator_in_y == tmp1179;
    assign tmp1183 = my_calculator_in_y == tmp8076;
    assign tmp1184 = tmp1180 | tmp1183;
    assign tmp1187 = my_calculator_in_y == tmp8080;
    assign tmp1188 = tmp1184 | tmp1187;
    assign tmp1189 = {tmp11[14], tmp11[13], tmp11[12], tmp11[11], tmp11[10], tmp11[9], tmp11[8], tmp11[7], tmp11[6], tmp11[5], tmp11[4], tmp11[3], tmp11[2], tmp11[1], tmp11[0]};
    assign tmp1195 = tmp2887 - tmp11;
    assign tmp1196 = {tmp1195[16]};
    assign tmp1202 = tmp150 ^ tmp152;
    assign tmp1208 = {tmp158[16]};
    assign tmp1214 = tmp162 ^ tmp6605;
    assign tmp1221 = {tmp579[16]};
    assign tmp1233 = {tmp183[16]};
    assign tmp1236 = tmp1233 ^ tmp6605;
    assign tmp1240 = tmp2887 == tmp141;
    assign tmp1258 = {tmp13[14], tmp13[13], tmp13[12], tmp13[11], tmp13[10], tmp13[9], tmp13[8], tmp13[7], tmp13[6], tmp13[5], tmp13[4], tmp13[3], tmp13[2], tmp13[1], tmp13[0]};
    assign tmp1259 = {tmp1258, const_135_0};
    assign tmp1265 = {tmp7254[16]};
    assign tmp1268 = tmp1265 ^ tmp6605;
    assign tmp1276 = tmp1259 - tmp2887;
    assign tmp1277 = {tmp1276[16]};
    assign tmp1280 = tmp1277 ^ tmp1307;
    assign tmp1283 = tmp1280 ^ tmp6605;
    assign tmp1284 = tmp558 & tmp1283;
    assign tmp1301 = tmp2887 - tmp1259;
    assign tmp1302 = {tmp1301[16]};
    assign tmp1305 = tmp1302 ^ tmp6605;
    assign tmp1306 = {tmp1259[15]};
    assign tmp1307 = ~tmp1306;
    assign tmp1308 = tmp1305 ^ tmp1307;
    assign tmp1309 = tmp2887 == tmp1259;
    assign tmp1310 = tmp1308 | tmp1309;
    assign tmp1311 = tmp7250 & tmp1310;
    assign tmp1312 = tmp1284 ? const_140_32767 : tmp1259;
    assign tmp1313 = tmp1311 ? _ver_out_tmp_55 : tmp1312;
    assign tmp1328 = {tmp274, const_142_0};
    assign tmp1340 = tmp1866 ^ tmp1905;
    assign tmp1347 = {tmp1328[15]};
    assign tmp1352 = tmp7511 ^ tmp6605;
    assign tmp1370 = tmp2887 - tmp1328;
    assign tmp1377 = tmp321 ^ tmp7538;
    assign tmp1379 = tmp1377 | tmp325;
    assign tmp1380 = tmp7154 & tmp1379;
    assign tmp1381 = tmp7515 ? const_147_32767 : tmp1328;
    assign tmp1397 = {tmp7641, const_149_0};
    assign tmp1403 = {tmp7280[16]};
    assign tmp1414 = tmp1397 - tmp2887;
    assign tmp1416 = {tmp1397[15]};
    assign tmp1418 = tmp7660 ^ tmp1445;
    assign tmp1422 = tmp7654 & tmp7666;
    assign tmp1429 = {tmp17[15]};
    assign tmp1440 = {tmp7684[16]};
    assign tmp1445 = ~tmp1416;
    assign tmp1446 = tmp7688 ^ tmp1445;
    assign tmp1448 = tmp1446 | tmp7692;
    assign tmp1449 = tmp2034 & tmp1448;
    assign tmp1451 = tmp1449 ? _ver_out_tmp_20 : tmp7695;
    assign tmp1464 = tmp1701 & tmp1188;
    assign tmp1467 = my_calculator_in_y == tmp8104;
    assign tmp1470 = my_calculator_in_y == tmp8108;
    assign tmp1471 = tmp1467 | tmp1470;
    assign tmp1484 = ~tmp1188;
    assign tmp1542 = ~tmp1133;
    assign tmp1555 = ~tmp1132;
    assign tmp1561 = tmp2078 & tmp1471;
    assign tmp1594 = my_calculator_in_y == tmp520;
    assign tmp1597 = my_calculator_in_y == tmp523;
    assign tmp1598 = tmp1594 | tmp1597;
    assign tmp1601 = {tmp2625, tmp11};
    assign tmp1604 = {tmp1629, tmp12};
    assign tmp1605 = tmp1601 + tmp1604;
    assign tmp1606 = {tmp1605[16], tmp1605[15], tmp1605[14], tmp1605[13], tmp1605[12], tmp1605[11], tmp1605[10], tmp1605[9], tmp1605[8], tmp1605[7], tmp1605[6], tmp1605[5], tmp1605[4], tmp1605[3], tmp1605[2], tmp1605[1], tmp1605[0]};
    assign tmp1607 = {tmp1606[15], tmp1606[14], tmp1606[13], tmp1606[12], tmp1606[11], tmp1606[10], tmp1606[9], tmp1606[8], tmp1606[7], tmp1606[6], tmp1606[5], tmp1606[4], tmp1606[3], tmp1606[2], tmp1606[1], tmp1606[0]};
    assign tmp1624 = tmp2887 - tmp12;
    assign tmp1625 = {tmp1624[16]};
    assign tmp1629 = {tmp12[15]};
    assign tmp1632 = tmp1202 & tmp667;
    assign tmp1637 = tmp1607 - tmp2887;
    assign tmp1638 = {tmp1637[16]};
    assign tmp1639 = {tmp1607[15]};
    assign tmp1640 = ~tmp1639;
    assign tmp1641 = tmp1638 ^ tmp1640;
    assign tmp1644 = tmp1641 ^ tmp6605;
    assign tmp1645 = tmp1607 == tmp2887;
    assign tmp1646 = tmp1644 | tmp1645;
    assign tmp1647 = tmp1632 & tmp1646;
    assign tmp1665 = {tmp2240[16]};
    assign tmp1672 = tmp586 & tmp2247;
    assign tmp1677 = tmp2887 - tmp1607;
    assign tmp1678 = {tmp1677[16]};
    assign tmp1681 = tmp1678 ^ tmp6605;
    assign tmp1684 = tmp1681 ^ tmp1640;
    assign tmp1686 = tmp1684 | tmp1645;
    assign tmp1687 = tmp1672 & tmp1686;
    assign tmp1688 = tmp1647 ? const_170_32767 : tmp1607;
    assign tmp1689 = tmp1687 ? _ver_out_tmp_61 : tmp1688;
    assign tmp1701 = tmp1841 & tmp1542;
    assign tmp1726 = {tmp593, tmp13};
    assign tmp1729 = {tmp650, tmp14};
    assign tmp1730 = tmp1726 + tmp1729;
    assign tmp1731 = {tmp1730[16], tmp1730[15], tmp1730[14], tmp1730[13], tmp1730[12], tmp1730[11], tmp1730[10], tmp1730[9], tmp1730[8], tmp1730[7], tmp1730[6], tmp1730[5], tmp1730[4], tmp1730[3], tmp1730[2], tmp1730[1], tmp1730[0]};
    assign tmp1732 = {tmp1731[15], tmp1731[14], tmp1731[13], tmp1731[12], tmp1731[11], tmp1731[10], tmp1731[9], tmp1731[8], tmp1731[7], tmp1731[6], tmp1731[5], tmp1731[4], tmp1731[3], tmp1731[2], tmp1731[1], tmp1731[0]};
    assign tmp1743 = ~tmp593;
    assign tmp1750 = {tmp2527[16]};
    assign tmp1753 = tmp1750 ^ tmp6605;
    assign tmp1757 = tmp558 & tmp679;
    assign tmp1762 = tmp1732 - tmp2887;
    assign tmp1763 = {tmp1762[16]};
    assign tmp1764 = {tmp1732[15]};
    assign tmp1765 = ~tmp1764;
    assign tmp1766 = tmp1763 ^ tmp1765;
    assign tmp1769 = tmp1766 ^ tmp6605;
    assign tmp1770 = tmp1732 == tmp2887;
    assign tmp1771 = tmp1769 | tmp1770;
    assign tmp1772 = tmp1757 & tmp1771;
    assign tmp1789 = tmp14 - tmp2887;
    assign tmp1790 = {tmp1789[16]};
    assign tmp1797 = tmp7250 & tmp6913;
    assign tmp1802 = tmp2887 - tmp1732;
    assign tmp1803 = {tmp1802[16]};
    assign tmp1806 = tmp1803 ^ tmp6605;
    assign tmp1809 = tmp1806 ^ tmp1765;
    assign tmp1811 = tmp1809 | tmp1770;
    assign tmp1812 = tmp1797 & tmp1811;
    assign tmp1813 = tmp1772 ? const_178_32767 : tmp1732;
    assign tmp1814 = tmp1812 ? _ver_out_tmp_59 : tmp1813;
    assign tmp1841 = tmp1141 & tmp1555;
    assign tmp1846 = ~tmp1471;
    assign tmp1849 = {tmp15[15]};
    assign tmp1854 = {tmp889, tmp16};
    assign tmp1855 = tmp770 + tmp1854;
    assign tmp1856 = {tmp1855[16], tmp1855[15], tmp1855[14], tmp1855[13], tmp1855[12], tmp1855[11], tmp1855[10], tmp1855[9], tmp1855[8], tmp1855[7], tmp1855[6], tmp1855[5], tmp1855[4], tmp1855[3], tmp1855[2], tmp1855[1], tmp1855[0]};
    assign tmp1857 = {tmp1856[15], tmp1856[14], tmp1856[13], tmp1856[12], tmp1856[11], tmp1856[10], tmp1856[9], tmp1856[8], tmp1856[7], tmp1856[6], tmp1856[5], tmp1856[4], tmp1856[3], tmp1856[2], tmp1856[1], tmp1856[0]};
    assign tmp1866 = tmp782 ^ tmp6605;
    assign tmp1882 = tmp1340 & tmp354;
    assign tmp1887 = tmp1857 - tmp2887;
    assign tmp1888 = {tmp1887[16]};
    assign tmp1889 = {tmp1857[15]};
    assign tmp1891 = tmp1888 ^ tmp1933;
    assign tmp1894 = tmp1891 ^ tmp6605;
    assign tmp1896 = tmp1894 | tmp1935;
    assign tmp1897 = tmp1882 & tmp1896;
    assign tmp1905 = ~tmp1849;
    assign tmp1922 = tmp7154 & tmp6825;
    assign tmp1927 = tmp2887 - tmp1857;
    assign tmp1928 = {tmp1927[16]};
    assign tmp1931 = tmp1928 ^ tmp6605;
    assign tmp1933 = ~tmp1889;
    assign tmp1934 = tmp1931 ^ tmp1933;
    assign tmp1935 = tmp2887 == tmp1857;
    assign tmp1936 = tmp1934 | tmp1935;
    assign tmp1937 = tmp1922 & tmp1936;
    assign tmp1938 = tmp1897 ? const_186_32767 : tmp1857;
    assign tmp1939 = tmp1937 ? _ver_out_tmp_64 : tmp1938;
    assign tmp1976 = {tmp1429, tmp17};
    assign tmp1979 = {tmp2041, tmp18};
    assign tmp1980 = tmp1976 + tmp1979;
    assign tmp1981 = {tmp1980[16], tmp1980[15], tmp1980[14], tmp1980[13], tmp1980[12], tmp1980[11], tmp1980[10], tmp1980[9], tmp1980[8], tmp1980[7], tmp1980[6], tmp1980[5], tmp1980[4], tmp1980[3], tmp1980[2], tmp1980[1], tmp1980[0]};
    assign tmp1982 = {tmp1981[15], tmp1981[14], tmp1981[13], tmp1981[12], tmp1981[11], tmp1981[10], tmp1981[9], tmp1981[8], tmp1981[7], tmp1981[6], tmp1981[5], tmp1981[4], tmp1981[3], tmp1981[2], tmp1981[1], tmp1981[0]};
    assign tmp1999 = tmp2887 - tmp18;
    assign tmp2006 = tmp918 ^ tmp6931;
    assign tmp2007 = tmp7654 & tmp2006;
    assign tmp2012 = tmp1982 - tmp2887;
    assign tmp2013 = {tmp2012[16]};
    assign tmp2015 = ~tmp2057;
    assign tmp2016 = tmp2013 ^ tmp2015;
    assign tmp2019 = tmp2016 ^ tmp6605;
    assign tmp2020 = tmp1982 == tmp2887;
    assign tmp2021 = tmp2019 | tmp2020;
    assign tmp2022 = tmp2007 & tmp2021;
    assign tmp2034 = tmp2343 ^ tmp6605;
    assign tmp2041 = {tmp18[15]};
    assign tmp2047 = tmp2034 & tmp6935;
    assign tmp2052 = tmp2887 - tmp1982;
    assign tmp2053 = {tmp2052[16]};
    assign tmp2056 = tmp2053 ^ tmp6605;
    assign tmp2057 = {tmp1982[15]};
    assign tmp2059 = tmp2056 ^ tmp2015;
    assign tmp2061 = tmp2059 | tmp2020;
    assign tmp2062 = tmp2047 & tmp2061;
    assign tmp2063 = tmp2022 ? const_194_32767 : tmp1982;
    assign tmp2064 = tmp2062 ? _ver_out_tmp_65 : tmp2063;
    assign tmp2078 = tmp1701 & tmp1484;
    assign tmp2081 = tmp2150 & tmp1598;
    assign tmp2099 = my_calculator_in_y == const_196_8;
    assign tmp2100 = tmp11 == _ver_out_tmp_87;
    assign tmp2106 = tmp2100 ? tmp6864 : tmp1195;
    assign tmp2125 = tmp2150 & tmp2151;
    assign tmp2126 = tmp2125 & tmp2099;
    assign tmp2150 = tmp2078 & tmp1846;
    assign tmp2151 = ~tmp1598;
    assign tmp2209 = {const_218_0, const_217_3};
    assign tmp2235 = tmp586 == tmp2247;
    assign tmp2240 = tmp12 - tmp2887;
    assign tmp2247 = tmp7186 ^ tmp6605;
    assign tmp2260 = tmp2247 == tmp7250;
    assign tmp2261 = tmp2235 & tmp2260;
    assign tmp2281 = ~tmp650;
    assign tmp2286 = tmp7250 == tmp6913;
    assign tmp2287 = tmp2261 & tmp2286;
    assign tmp2322 = tmp7154 == tmp6825;
    assign tmp2343 = tmp834 ^ tmp7675;
    assign tmp2347 = tmp6825 == tmp2034;
    assign tmp2348 = tmp2322 & tmp2347;
    assign tmp2353 = tmp17 - tmp2887;
    assign tmp2365 = tmp18 - tmp2887;
    assign tmp2366 = {tmp2365[16]};
    assign tmp2369 = tmp2366 ^ tmp6931;
    assign tmp2373 = tmp2034 == tmp6935;
    assign tmp2374 = tmp2348 & tmp2373;
    assign tmp2387 = tmp15 == tmp2887;
    assign tmp2390 = tmp16 == tmp2887;
    assign tmp2391 = tmp2387 | tmp2390;
    assign tmp2395 = tmp2391 | tmp2759;
    assign tmp2398 = tmp18 == tmp2887;
    assign tmp2399 = tmp2395 | tmp2398;
    assign tmp2410 = tmp8034 & tmp8035;
    assign tmp2411 = ~tmp8036;
    assign tmp2412 = tmp2410 & tmp2411;
    assign tmp2423 = {tmp11[0]};
    assign tmp2424 = {tmp12[0]};
    assign tmp2425 = tmp2423 | tmp2424;
    assign tmp2426 = {tmp13[0]};
    assign tmp2427 = tmp2425 | tmp2426;
    assign tmp2428 = {tmp14[0]};
    assign tmp2429 = tmp2427 | tmp2428;
    assign tmp2430 = ~tmp2429;
    assign tmp2453 = tmp8037 & tmp586;
    assign tmp2458 = tmp15 - tmp2887;
    assign tmp2466 = tmp2453 & tmp7154;
    assign tmp2474 = {tmp2106[15], tmp2106[14], tmp2106[13], tmp2106[12], tmp2106[11], tmp2106[10], tmp2106[9], tmp2106[8], tmp2106[7], tmp2106[6], tmp2106[5], tmp2106[4], tmp2106[3], tmp2106[2], tmp2106[1], tmp2106[0]};
    assign tmp2486 = tmp12 == _ver_out_tmp_82;
    assign tmp2492 = tmp2486 ? tmp6864 : tmp1624;
    assign tmp2512 = {tmp6865[15], tmp6865[14], tmp6865[13], tmp6865[12], tmp6865[11], tmp6865[10], tmp6865[9], tmp6865[8], tmp6865[7], tmp6865[6], tmp6865[5], tmp6865[4], tmp6865[3], tmp6865[2], tmp6865[1], tmp6865[0]};
    assign tmp2524 = tmp14 == _ver_out_tmp_86;
    assign tmp2527 = tmp2887 - tmp14;
    assign tmp2530 = tmp2524 ? tmp6864 : tmp2527;
    assign tmp2531 = {tmp2530[15], tmp2530[14], tmp2530[13], tmp2530[12], tmp2530[11], tmp2530[10], tmp2530[9], tmp2530[8], tmp2530[7], tmp2530[6], tmp2530[5], tmp2530[4], tmp2530[3], tmp2530[2], tmp2530[1], tmp2530[0]};
    assign tmp2549 = tmp6772 ? tmp6864 : tmp7495;
    assign tmp2550 = {tmp2549[15], tmp2549[14], tmp2549[13], tmp2549[12], tmp2549[11], tmp2549[10], tmp2549[9], tmp2549[8], tmp2549[7], tmp2549[6], tmp2549[5], tmp2549[4], tmp2549[3], tmp2549[2], tmp2549[1], tmp2549[0]};
    assign tmp2561 = tmp2681 & tmp2466;
    assign tmp2565 = tmp2887 - tmp16;
    assign tmp2569 = {tmp1092[15], tmp1092[14], tmp1092[13], tmp1092[12], tmp1092[11], tmp1092[10], tmp1092[9], tmp1092[8], tmp1092[7], tmp1092[6], tmp1092[5], tmp1092[4], tmp1092[3], tmp1092[2], tmp1092[1], tmp1092[0]};
    assign tmp2581 = tmp17 == _ver_out_tmp_0;
    assign tmp2588 = {tmp6887[15], tmp6887[14], tmp6887[13], tmp6887[12], tmp6887[11], tmp6887[10], tmp6887[9], tmp6887[8], tmp6887[7], tmp6887[6], tmp6887[5], tmp6887[4], tmp6887[3], tmp6887[2], tmp6887[1], tmp6887[0]};
    assign tmp2606 = tmp6936 ? tmp6864 : tmp1999;
    assign tmp2607 = {tmp2606[15], tmp2606[14], tmp2606[13], tmp2606[12], tmp2606[11], tmp2606[10], tmp2606[9], tmp2606[8], tmp2606[7], tmp2606[6], tmp2606[5], tmp2606[4], tmp2606[3], tmp2606[2], tmp2606[1], tmp2606[0]};
    assign tmp2610 = tmp2646 & tmp4395;
    assign tmp2625 = {tmp11[15]};
    assign tmp2627 = tmp1221 ^ tmp152;
    assign tmp2643 = tmp586 & tmp7154;
    assign tmp2644 = ~tmp2643;
    assign tmp2645 = tmp8037 & tmp2644;
    assign tmp2646 = ~tmp33;
    assign tmp2649 = ~tmp37;
    assign tmp2681 = tmp4999 & tmp8129;
    assign tmp2722 = tmp2681 & tmp2747;
    assign tmp2736 = tmp2722 & tmp2645;
    assign tmp2747 = ~tmp2466;
    assign tmp2756 = tmp2387 & tmp2390;
    assign tmp2759 = tmp17 == tmp2887;
    assign tmp2760 = tmp2756 & tmp2759;
    assign tmp2764 = tmp2760 & tmp2398;
    assign tmp2775 = tmp2681 & tmp2764;
    assign tmp2807 = tmp6765 ^ tmp1905;
    assign tmp2811 = tmp586 == tmp7154;
    assign tmp2812 = ~tmp2811;
    assign tmp2826 = tmp6183 & tmp2812;
    assign tmp2870 = {tmp2492[15], tmp2492[14], tmp2492[13], tmp2492[12], tmp2492[11], tmp2492[10], tmp2492[9], tmp2492[8], tmp2492[7], tmp2492[6], tmp2492[5], tmp2492[4], tmp2492[3], tmp2492[2], tmp2492[1], tmp2492[0]};
    assign tmp2885 = tmp13 == _ver_out_tmp_9;
    assign tmp2887 = {tmp143, const_308_0};
    assign tmp2935 = tmp8058 - tmp3602;
    assign tmp2936 = {tmp2935[16]};
    assign tmp2937 = {tmp3602[15]};
    assign tmp2939 = tmp2936 ^ tmp3608;
    assign tmp2942 = tmp2939 ^ tmp5173;
    assign tmp2943 = tmp3602 == tmp8058;
    assign tmp2944 = tmp2942 | tmp2943;
    assign tmp2948 = {tmp4860, tmp3614};
    assign tmp2951 = tmp8062 - tmp2948;
    assign tmp2952 = {tmp2951[16]};
    assign tmp2953 = {tmp2948[15]};
    assign tmp2954 = ~tmp2953;
    assign tmp2955 = tmp2952 ^ tmp2954;
    assign tmp2958 = tmp2955 ^ tmp3360;
    assign tmp2959 = tmp2948 == tmp8062;
    assign tmp2960 = tmp2958 | tmp2959;
    assign tmp2961 = tmp2944 & tmp2960;
    assign tmp2968 = tmp8066 - tmp4890;
    assign tmp2969 = {tmp2968[16]};
    assign tmp2970 = {tmp4890[15]};
    assign tmp2972 = tmp2969 ^ tmp3638;
    assign tmp2975 = tmp2972 ^ tmp4652;
    assign tmp2976 = tmp4890 == tmp8066;
    assign tmp2977 = tmp2975 | tmp2976;
    assign tmp2978 = tmp2961 & tmp2977;
    assign tmp2982 = {tmp4916, tmp4915};
    assign tmp2985 = tmp8070 - tmp2982;
    assign tmp2986 = {tmp2985[16]};
    assign tmp2987 = {tmp2982[15]};
    assign tmp2988 = ~tmp2987;
    assign tmp2989 = tmp2986 ^ tmp2988;
    assign tmp2992 = tmp2989 ^ tmp3486;
    assign tmp2993 = tmp2982 == tmp8070;
    assign tmp2994 = tmp2992 | tmp2993;
    assign tmp2995 = tmp2978 & tmp2994;
    assign tmp3029 = {tmp3599[14]};
    assign tmp3145 = tmp3397 & tmp8038;
    assign tmp3196 = ~tmp8038;
    assign tmp3215 = tmp3397 & tmp3196;
    assign tmp3253 = {tmp5139, const_319_0};
    assign tmp3263 = {tmp8058[15]};
    assign tmp3270 = tmp3253 - tmp2887;
    assign tmp3271 = {tmp3270[16]};
    assign tmp3274 = tmp3271 ^ tmp5550;
    assign tmp3278 = tmp4497 & tmp5164;
    assign tmp3284 = {tmp5170[16]};
    assign tmp3287 = tmp3284 ^ tmp5173;
    assign tmp3290 = tmp3287 ^ tmp6605;
    assign tmp3307 = tmp5192 ? _ver_out_tmp_15 : tmp5193;
    assign tmp3327 = {tmp5663, const_326_0};
    assign tmp3345 = {tmp5681[16]};
    assign tmp3347 = ~tmp5683;
    assign tmp3348 = tmp3345 ^ tmp3347;
    assign tmp3351 = tmp3348 ^ tmp6605;
    assign tmp3360 = ~tmp4573;
    assign tmp3361 = tmp4594 ^ tmp3360;
    assign tmp3373 = tmp5707 ^ tmp6605;
    assign tmp3376 = tmp3373 ^ tmp3347;
    assign tmp3379 = tmp5701 & tmp5272;
    assign tmp3397 = tmp5209 & tmp2995;
    assign tmp3413 = tmp5311 ^ tmp4652;
    assign tmp3419 = {tmp5815[16]};
    assign tmp3435 = tmp5829 ^ tmp4652;
    assign tmp3453 = tmp5835 & tmp5353;
    assign tmp3480 = tmp2887 - tmp8070;
    assign tmp3486 = ~tmp4729;
    assign tmp3496 = tmp5401 ^ tmp5952;
    assign tmp3506 = {tmp5962[16]};
    assign tmp3521 = tmp5426 ^ tmp6605;
    assign tmp3526 = tmp5432 | tmp5982;
    assign tmp3528 = tmp5957 ? const_345_32767 : tmp5932;
    assign tmp3550 = tmp8058 - tmp8042;
    assign tmp3553 = ~tmp4481;
    assign tmp3554 = tmp4477 ^ tmp3553;
    assign tmp3557 = tmp3554 ^ tmp5173;
    assign tmp3558 = tmp8042 == tmp8058;
    assign tmp3559 = tmp3557 | tmp3558;
    assign tmp3566 = tmp4554 ^ tmp4623;
    assign tmp3569 = tmp3566 ^ tmp3360;
    assign tmp3570 = tmp8046 == tmp8062;
    assign tmp3571 = tmp3569 | tmp3570;
    assign tmp3572 = tmp3559 & tmp3571;
    assign tmp3575 = tmp8066 - tmp8050;
    assign tmp3576 = {tmp3575[16]};
    assign tmp3579 = tmp3576 ^ tmp4257;
    assign tmp3582 = tmp3579 ^ tmp4652;
    assign tmp3583 = tmp8050 == tmp8066;
    assign tmp3584 = tmp3582 | tmp3583;
    assign tmp3585 = tmp3572 & tmp3584;
    assign tmp3588 = tmp8070 - tmp8054;
    assign tmp3589 = {tmp3588[16]};
    assign tmp3592 = tmp3589 ^ tmp6543;
    assign tmp3595 = tmp3592 ^ tmp3486;
    assign tmp3596 = tmp8054 == tmp8070;
    assign tmp3597 = tmp3595 | tmp3596;
    assign tmp3598 = tmp3585 & tmp3597;
    assign tmp3599 = {tmp8042[15], tmp8042[14], tmp8042[13], tmp8042[12], tmp8042[11], tmp8042[10], tmp8042[9], tmp8042[8], tmp8042[7], tmp8042[6], tmp8042[5], tmp8042[4], tmp8042[3], tmp8042[2], tmp8042[1]};
    assign tmp3602 = {tmp3029, tmp3599};
    assign tmp3605 = tmp3602 - tmp8058;
    assign tmp3606 = {tmp3605[16]};
    assign tmp3608 = ~tmp2937;
    assign tmp3609 = tmp3606 ^ tmp3608;
    assign tmp3612 = tmp3609 ^ tmp5173;
    assign tmp3613 = tmp3598 & tmp3612;
    assign tmp3614 = {tmp8046[15], tmp8046[14], tmp8046[13], tmp8046[12], tmp8046[11], tmp8046[10], tmp8046[9], tmp8046[8], tmp8046[7], tmp8046[6], tmp8046[5], tmp8046[4], tmp8046[3], tmp8046[2], tmp8046[1]};
    assign tmp3620 = tmp2948 - tmp8062;
    assign tmp3621 = {tmp3620[16]};
    assign tmp3624 = tmp3621 ^ tmp2954;
    assign tmp3627 = tmp3624 ^ tmp3360;
    assign tmp3628 = tmp3613 & tmp3627;
    assign tmp3630 = {tmp4887[14]};
    assign tmp3635 = tmp4890 - tmp8066;
    assign tmp3636 = {tmp3635[16]};
    assign tmp3638 = ~tmp2970;
    assign tmp3639 = tmp3636 ^ tmp3638;
    assign tmp3640 = {tmp8066[15]};
    assign tmp3642 = tmp3639 ^ tmp4652;
    assign tmp3643 = tmp3628 & tmp3642;
    assign tmp3650 = tmp2982 - tmp8070;
    assign tmp3651 = {tmp3650[16]};
    assign tmp3654 = tmp3651 ^ tmp2988;
    assign tmp3657 = tmp3654 ^ tmp3486;
    assign tmp3658 = tmp3643 & tmp3657;
    assign tmp3694 = tmp6656 & tmp3658;
    assign tmp3713 = _ver_out_tmp_27 == tmp8058;
    assign tmp3719 = tmp3713 ? tmp6864 : tmp5145;
    assign tmp3721 = {tmp4481, tmp4481};
    assign tmp3722 = {tmp3721, tmp8042};
    assign tmp3725 = {tmp6083, tmp3719};
    assign tmp3726 = tmp3722 + tmp3725;
    assign tmp3727 = {tmp3726[17], tmp3726[16], tmp3726[15], tmp3726[14], tmp3726[13], tmp3726[12], tmp3726[11], tmp3726[10], tmp3726[9], tmp3726[8], tmp3726[7], tmp3726[6], tmp3726[5], tmp3726[4], tmp3726[3], tmp3726[2], tmp3726[1], tmp3726[0]};
    assign tmp3728 = {tmp3727[15], tmp3727[14], tmp3727[13], tmp3727[12], tmp3727[11], tmp3727[10], tmp3727[9], tmp3727[8], tmp3727[7], tmp3727[6], tmp3727[5], tmp3727[4], tmp3727[3], tmp3727[2], tmp3727[1], tmp3727[0]};
    assign tmp3733 = tmp2887 - tmp8042;
    assign tmp3734 = {tmp3733[16]};
    assign tmp3737 = tmp3734 ^ tmp6605;
    assign tmp3742 = {const_355_0, const_355_0, const_355_0, const_355_0, const_355_0, const_355_0, const_355_0, const_355_0, const_355_0, const_355_0, const_355_0, const_355_0, const_355_0, const_355_0, const_355_0, const_355_0};
    assign tmp3745 = tmp6440 - tmp3719;
    assign tmp3746 = {tmp3745[17]};
    assign tmp3752 = tmp6109 ^ tmp3788;
    assign tmp3753 = tmp6100 & tmp3752;
    assign tmp3758 = tmp3728 - tmp2887;
    assign tmp3759 = {tmp3758[16]};
    assign tmp3760 = {tmp3728[15]};
    assign tmp3762 = tmp3759 ^ tmp6164;
    assign tmp3765 = tmp3762 ^ tmp6605;
    assign tmp3766 = tmp3728 == tmp2887;
    assign tmp3773 = tmp8042 - tmp2887;
    assign tmp3777 = tmp5495 ^ tmp3553;
    assign tmp3780 = tmp3777 ^ tmp6605;
    assign tmp3785 = tmp3719 - tmp6440;
    assign tmp3786 = {tmp3785[17]};
    assign tmp3788 = ~tmp6083;
    assign tmp3793 = tmp3780 & tmp6152;
    assign tmp3798 = tmp2887 - tmp3728;
    assign tmp3802 = tmp6159 ^ tmp6605;
    assign tmp3810 = tmp6168 ? _ver_out_tmp_31 : tmp6169;
    assign tmp3856 = {tmp6229, tmp8046};
    assign tmp3860 = tmp3856 + tmp6233;
    assign tmp3861 = {tmp3860[17], tmp3860[16], tmp3860[15], tmp3860[14], tmp3860[13], tmp3860[12], tmp3860[11], tmp3860[10], tmp3860[9], tmp3860[8], tmp3860[7], tmp3860[6], tmp3860[5], tmp3860[4], tmp3860[3], tmp3860[2], tmp3860[1], tmp3860[0]};
    assign tmp3867 = tmp2887 - tmp8046;
    assign tmp3880 = {tmp6253[17]};
    assign tmp3892 = tmp6236 - tmp2887;
    assign tmp3893 = {tmp3892[16]};
    assign tmp3901 = tmp6273 | tmp3940;
    assign tmp3919 = tmp6227 - tmp6440;
    assign tmp3921 = {tmp6227[16]};
    assign tmp3922 = ~tmp3921;
    assign tmp3926 = tmp6297 ^ tmp4016;
    assign tmp3937 = {tmp6236[15]};
    assign tmp3939 = tmp6310 ^ tmp6312;
    assign tmp3940 = tmp2887 == tmp6236;
    assign tmp3941 = tmp3939 | tmp3940;
    assign tmp3943 = tmp6276 ? const_373_32767 : tmp6236;
    assign tmp3944 = tmp6316 ? _ver_out_tmp_35 : tmp3943;
    assign tmp3987 = tmp6369 ? tmp6864 : tmp5803;
    assign tmp3988 = {tmp8050[15]};
    assign tmp3990 = {tmp6377, tmp8050};
    assign tmp3991 = {tmp3987[16]};
    assign tmp3995 = {tmp6382[17], tmp6382[16], tmp6382[15], tmp6382[14], tmp6382[13], tmp6382[12], tmp6382[11], tmp6382[10], tmp6382[9], tmp6382[8], tmp6382[7], tmp6382[6], tmp6382[5], tmp6382[4], tmp6382[3], tmp6382[2], tmp6382[1], tmp6382[0]};
    assign tmp3996 = {tmp3995[15], tmp3995[14], tmp3995[13], tmp3995[12], tmp3995[11], tmp3995[10], tmp3995[9], tmp3995[8], tmp3995[7], tmp3995[6], tmp3995[5], tmp3995[4], tmp3995[3], tmp3995[2], tmp3995[1], tmp3995[0]};
    assign tmp4001 = tmp2887 - tmp8050;
    assign tmp4008 = tmp5740 ^ tmp4257;
    assign tmp4013 = tmp6440 - tmp3987;
    assign tmp4014 = {tmp4013[17]};
    assign tmp4016 = ~tmp6107;
    assign tmp4017 = tmp4014 ^ tmp4016;
    assign tmp4021 = tmp4008 & tmp6408;
    assign tmp4026 = tmp3996 - tmp2887;
    assign tmp4027 = {tmp4026[16]};
    assign tmp4030 = tmp4027 ^ tmp4072;
    assign tmp4033 = tmp4030 ^ tmp6605;
    assign tmp4035 = tmp4033 | tmp6462;
    assign tmp4036 = tmp4021 & tmp4035;
    assign tmp4041 = tmp8050 - tmp2887;
    assign tmp4045 = tmp6430 ^ tmp4257;
    assign tmp4053 = tmp3987 - tmp6440;
    assign tmp4054 = {tmp4053[17]};
    assign tmp4056 = ~tmp3991;
    assign tmp4057 = tmp4054 ^ tmp4056;
    assign tmp4060 = tmp4057 ^ tmp4016;
    assign tmp4061 = tmp5768 & tmp4060;
    assign tmp4066 = tmp2887 - tmp3996;
    assign tmp4067 = {tmp4066[16]};
    assign tmp4070 = tmp4067 ^ tmp6605;
    assign tmp4071 = {tmp3996[15]};
    assign tmp4072 = ~tmp4071;
    assign tmp4073 = tmp4070 ^ tmp4072;
    assign tmp4076 = tmp4061 & tmp6463;
    assign tmp4077 = tmp4036 ? const_386_32767 : tmp3996;
    assign tmp4078 = tmp4076 ? _ver_out_tmp_41 : tmp4077;
    assign tmp4123 = {tmp6542, tmp6542};
    assign tmp4127 = {tmp6591, tmp6523};
    assign tmp4128 = tmp6526 + tmp4127;
    assign tmp4129 = {tmp4128[17], tmp4128[16], tmp4128[15], tmp4128[14], tmp4128[13], tmp4128[12], tmp4128[11], tmp4128[10], tmp4128[9], tmp4128[8], tmp4128[7], tmp4128[6], tmp4128[5], tmp4128[4], tmp4128[3], tmp4128[2], tmp4128[1], tmp4128[0]};
    assign tmp4130 = {tmp4129[15], tmp4129[14], tmp4129[13], tmp4129[12], tmp4129[11], tmp4129[10], tmp4129[9], tmp4129[8], tmp4129[7], tmp4129[6], tmp4129[5], tmp4129[4], tmp4129[3], tmp4129[2], tmp4129[1], tmp4129[0]};
    assign tmp4135 = tmp2887 - tmp8054;
    assign tmp4142 = tmp5874 ^ tmp6543;
    assign tmp4153 = ~tmp6591;
    assign tmp4155 = tmp4142 & tmp6556;
    assign tmp4168 = tmp4130 == tmp2887;
    assign tmp4169 = tmp6569 | tmp4168;
    assign tmp4170 = tmp4155 & tmp4169;
    assign tmp4182 = tmp5899 ^ tmp6605;
    assign tmp4187 = tmp6523 - tmp6440;
    assign tmp4207 = tmp6606 ^ tmp6608;
    assign tmp4209 = tmp4207 | tmp4168;
    assign tmp4210 = tmp6597 & tmp4209;
    assign tmp4212 = tmp4210 ? _ver_out_tmp_46 : tmp6613;
    assign tmp4233 = tmp8042 - tmp8058;
    assign tmp4234 = {tmp4233[16]};
    assign tmp4237 = tmp4234 ^ tmp3553;
    assign tmp4240 = tmp4237 ^ tmp5173;
    assign tmp4243 = tmp8046 - tmp8062;
    assign tmp4244 = {tmp4243[16]};
    assign tmp4247 = tmp4244 ^ tmp4623;
    assign tmp4250 = tmp4247 ^ tmp3360;
    assign tmp4251 = tmp4240 & tmp4250;
    assign tmp4254 = tmp8050 - tmp8066;
    assign tmp4255 = {tmp4254[16]};
    assign tmp4257 = ~tmp3988;
    assign tmp4258 = tmp4255 ^ tmp4257;
    assign tmp4261 = tmp4258 ^ tmp4652;
    assign tmp4262 = tmp4251 & tmp4261;
    assign tmp4265 = tmp8054 - tmp8070;
    assign tmp4266 = {tmp4265[16]};
    assign tmp4269 = tmp4266 ^ tmp6543;
    assign tmp4272 = tmp4269 ^ tmp3486;
    assign tmp4273 = tmp4262 & tmp4272;
    assign tmp4395 = ~tmp36;
    assign tmp4413 = tmp6633 & tmp4273;
    assign tmp4469 = ~tmp2995;
    assign tmp4477 = {tmp3550[16]};
    assign tmp4480 = tmp4477 ^ tmp5173;
    assign tmp4481 = {tmp8042[15]};
    assign tmp4483 = tmp4480 ^ tmp3553;
    assign tmp4484 = {tmp8058[13], tmp8058[12], tmp8058[11], tmp8058[10], tmp8058[9], tmp8058[8], tmp8058[7], tmp8058[6], tmp8058[5], tmp8058[4], tmp8058[3], tmp8058[2], tmp8058[1], tmp8058[0]};
    assign tmp4485 = {tmp4484, const_403_0};
    assign tmp4494 = tmp5146 ^ tmp6605;
    assign tmp4497 = tmp4494 ^ tmp5173;
    assign tmp4502 = tmp4485 - tmp2887;
    assign tmp4503 = {tmp4502[16]};
    assign tmp4504 = {tmp4485[15]};
    assign tmp4505 = ~tmp4504;
    assign tmp4506 = tmp4503 ^ tmp4505;
    assign tmp4509 = tmp4506 ^ tmp6605;
    assign tmp4510 = tmp4497 & tmp4509;
    assign tmp4527 = tmp2887 - tmp4485;
    assign tmp4528 = {tmp4527[16]};
    assign tmp4531 = tmp4528 ^ tmp6605;
    assign tmp4534 = tmp4531 ^ tmp4505;
    assign tmp4535 = tmp2887 == tmp4485;
    assign tmp4536 = tmp4534 | tmp4535;
    assign tmp4537 = tmp3290 & tmp4536;
    assign tmp4538 = tmp4510 ? const_408_32767 : tmp4485;
    assign tmp4539 = tmp4537 ? _ver_out_tmp_49 : tmp4538;
    assign tmp4542 = tmp8042 - tmp4539;
    assign tmp4543 = {tmp4542[16]};
    assign tmp4546 = tmp4543 ^ tmp3553;
    assign tmp4547 = {tmp4539[15]};
    assign tmp4548 = ~tmp4547;
    assign tmp4549 = tmp4546 ^ tmp4548;
    assign tmp4550 = tmp4483 & tmp4549;
    assign tmp4553 = tmp8062 - tmp8046;
    assign tmp4554 = {tmp4553[16]};
    assign tmp4557 = tmp4554 ^ tmp3360;
    assign tmp4560 = tmp4557 ^ tmp4623;
    assign tmp4561 = tmp4550 & tmp4560;
    assign tmp4562 = {tmp8062[13], tmp8062[12], tmp8062[11], tmp8062[10], tmp8062[9], tmp8062[8], tmp8062[7], tmp8062[6], tmp8062[5], tmp8062[4], tmp8062[3], tmp8062[2], tmp8062[1], tmp8062[0]};
    assign tmp4563 = {tmp4562, const_410_0};
    assign tmp4573 = {tmp8062[15]};
    assign tmp4575 = tmp5673 ^ tmp3360;
    assign tmp4580 = tmp4563 - tmp2887;
    assign tmp4581 = {tmp4580[16]};
    assign tmp4582 = {tmp4563[15]};
    assign tmp4583 = ~tmp4582;
    assign tmp4584 = tmp4581 ^ tmp4583;
    assign tmp4587 = tmp4584 ^ tmp6605;
    assign tmp4588 = tmp4575 & tmp4587;
    assign tmp4594 = {tmp5694[16]};
    assign tmp4605 = tmp2887 - tmp4563;
    assign tmp4606 = {tmp4605[16]};
    assign tmp4609 = tmp4606 ^ tmp6605;
    assign tmp4612 = tmp4609 ^ tmp4583;
    assign tmp4613 = tmp2887 == tmp4563;
    assign tmp4614 = tmp4612 | tmp4613;
    assign tmp4615 = tmp5701 & tmp4614;
    assign tmp4616 = tmp4588 ? const_415_32767 : tmp4563;
    assign tmp4617 = tmp4615 ? _ver_out_tmp_50 : tmp4616;
    assign tmp4620 = tmp8046 - tmp4617;
    assign tmp4621 = {tmp4620[16]};
    assign tmp4623 = ~tmp5607;
    assign tmp4624 = tmp4621 ^ tmp4623;
    assign tmp4625 = {tmp4617[15]};
    assign tmp4626 = ~tmp4625;
    assign tmp4627 = tmp4624 ^ tmp4626;
    assign tmp4628 = tmp4561 & tmp4627;
    assign tmp4635 = tmp3576 ^ tmp4652;
    assign tmp4638 = tmp4635 ^ tmp4257;
    assign tmp4639 = tmp4628 & tmp4638;
    assign tmp4640 = {tmp8066[13], tmp8066[12], tmp8066[11], tmp8066[10], tmp8066[9], tmp8066[8], tmp8066[7], tmp8066[6], tmp8066[5], tmp8066[4], tmp8066[3], tmp8066[2], tmp8066[1], tmp8066[0]};
    assign tmp4641 = {tmp4640, const_417_0};
    assign tmp4652 = ~tmp3640;
    assign tmp4658 = tmp4641 - tmp2887;
    assign tmp4659 = {tmp4658[16]};
    assign tmp4660 = {tmp4641[15]};
    assign tmp4661 = ~tmp4660;
    assign tmp4662 = tmp4659 ^ tmp4661;
    assign tmp4665 = tmp4662 ^ tmp6605;
    assign tmp4666 = tmp3413 & tmp4665;
    assign tmp4683 = tmp2887 - tmp4641;
    assign tmp4684 = {tmp4683[16]};
    assign tmp4687 = tmp4684 ^ tmp6605;
    assign tmp4690 = tmp4687 ^ tmp4661;
    assign tmp4691 = tmp2887 == tmp4641;
    assign tmp4692 = tmp4690 | tmp4691;
    assign tmp4693 = tmp5835 & tmp4692;
    assign tmp4694 = tmp4666 ? const_422_32767 : tmp4641;
    assign tmp4695 = tmp4693 ? _ver_out_tmp_51 : tmp4694;
    assign tmp4698 = tmp8050 - tmp4695;
    assign tmp4699 = {tmp4698[16]};
    assign tmp4702 = tmp4699 ^ tmp4257;
    assign tmp4703 = {tmp4695[15]};
    assign tmp4704 = ~tmp4703;
    assign tmp4705 = tmp4702 ^ tmp4704;
    assign tmp4706 = tmp4639 & tmp4705;
    assign tmp4713 = tmp3589 ^ tmp3486;
    assign tmp4716 = tmp4713 ^ tmp6543;
    assign tmp4717 = tmp4706 & tmp4716;
    assign tmp4718 = {tmp8070[13], tmp8070[12], tmp8070[11], tmp8070[10], tmp8070[9], tmp8070[8], tmp8070[7], tmp8070[6], tmp8070[5], tmp8070[4], tmp8070[3], tmp8070[2], tmp8070[1], tmp8070[0]};
    assign tmp4719 = {tmp4718, const_424_0};
    assign tmp4725 = {tmp3480[16]};
    assign tmp4729 = {tmp8070[15]};
    assign tmp4736 = tmp4719 - tmp2887;
    assign tmp4737 = {tmp4736[16]};
    assign tmp4740 = tmp4737 ^ tmp4767;
    assign tmp4743 = tmp4740 ^ tmp6605;
    assign tmp4744 = tmp5395 & tmp4743;
    assign tmp4761 = tmp2887 - tmp4719;
    assign tmp4762 = {tmp4761[16]};
    assign tmp4765 = tmp4762 ^ tmp6605;
    assign tmp4766 = {tmp4719[15]};
    assign tmp4767 = ~tmp4766;
    assign tmp4768 = tmp4765 ^ tmp4767;
    assign tmp4769 = tmp2887 == tmp4719;
    assign tmp4770 = tmp4768 | tmp4769;
    assign tmp4771 = tmp5420 & tmp4770;
    assign tmp4772 = tmp4744 ? const_429_32767 : tmp4719;
    assign tmp4773 = tmp4771 ? _ver_out_tmp_54 : tmp4772;
    assign tmp4776 = tmp8054 - tmp4773;
    assign tmp4777 = {tmp4776[16]};
    assign tmp4780 = tmp4777 ^ tmp6543;
    assign tmp4781 = {tmp4773[15]};
    assign tmp4782 = ~tmp4781;
    assign tmp4783 = tmp4780 ^ tmp4782;
    assign tmp4784 = tmp4717 & tmp4783;
    assign tmp4860 = {tmp3614[14]};
    assign tmp4886 = tmp5013 & tmp8038;
    assign tmp4887 = {tmp8050[15], tmp8050[14], tmp8050[13], tmp8050[12], tmp8050[11], tmp8050[10], tmp8050[9], tmp8050[8], tmp8050[7], tmp8050[6], tmp8050[5], tmp8050[4], tmp8050[3], tmp8050[2], tmp8050[1]};
    assign tmp4890 = {tmp3630, tmp4887};
    assign tmp4915 = {tmp8054[15], tmp8054[14], tmp8054[13], tmp8054[12], tmp8054[11], tmp8054[10], tmp8054[9], tmp8054[8], tmp8054[7], tmp8054[6], tmp8054[5], tmp8054[4], tmp8054[3], tmp8054[2], tmp8054[1]};
    assign tmp4916 = {tmp4915[14]};
    assign tmp4971 = tmp2610 & tmp2649;
    assign tmp4999 = tmp7818 & tmp7628;
    assign tmp5011 = tmp6633 & tmp6634;
    assign tmp5013 = tmp5011 & tmp4784;
    assign tmp5102 = ~tmp2812;
    assign tmp5139 = {tmp8058[14], tmp8058[13], tmp8058[12], tmp8058[11], tmp8058[10], tmp8058[9], tmp8058[8], tmp8058[7], tmp8058[6], tmp8058[5], tmp8058[4], tmp8058[3], tmp8058[2], tmp8058[1], tmp8058[0]};
    assign tmp5145 = tmp2887 - tmp8058;
    assign tmp5146 = {tmp5145[16]};
    assign tmp5164 = tmp3274 ^ tmp6605;
    assign tmp5170 = tmp8058 - tmp2887;
    assign tmp5173 = ~tmp3263;
    assign tmp5182 = tmp2887 - tmp3253;
    assign tmp5187 = {tmp3253[15]};
    assign tmp5189 = tmp5576 ^ tmp5550;
    assign tmp5192 = tmp3290 & tmp5581;
    assign tmp5193 = tmp3278 ? const_438_32767 : tmp3253;
    assign tmp5209 = tmp6183 & tmp5102;
    assign tmp5219 = tmp5013 & tmp3196;
    assign tmp5271 = tmp2887 == tmp3327;
    assign tmp5272 = tmp3376 | tmp5271;
    assign tmp5274 = tmp5689 ? const_445_32767 : tmp3327;
    assign tmp5301 = {tmp8066[14], tmp8066[13], tmp8066[12], tmp8066[11], tmp8066[10], tmp8066[9], tmp8066[8], tmp8066[7], tmp8066[6], tmp8066[5], tmp8066[4], tmp8066[3], tmp8066[2], tmp8066[1], tmp8066[0]};
    assign tmp5311 = tmp5804 ^ tmp6605;
    assign tmp5323 = tmp3419 ^ tmp5846;
    assign tmp5326 = tmp5323 ^ tmp6605;
    assign tmp5327 = tmp3413 & tmp5326;
    assign tmp5345 = {tmp5840[16]};
    assign tmp5352 = tmp2887 == tmp5798;
    assign tmp5353 = tmp5847 | tmp5352;
    assign tmp5356 = tmp3453 ? _ver_out_tmp_58 : tmp5851;
    assign tmp5395 = tmp5941 ^ tmp3486;
    assign tmp5400 = tmp5932 - tmp2887;
    assign tmp5401 = {tmp5400[16]};
    assign tmp5402 = {tmp5932[15]};
    assign tmp5417 = tmp3506 ^ tmp3486;
    assign tmp5420 = tmp5417 ^ tmp6605;
    assign tmp5425 = tmp2887 - tmp5932;
    assign tmp5426 = {tmp5425[16]};
    assign tmp5432 = tmp3521 ^ tmp5952;
    assign tmp5435 = tmp5420 & tmp3526;
    assign tmp5463 = {tmp8042[14], tmp8042[13], tmp8042[12], tmp8042[11], tmp8042[10], tmp8042[9], tmp8042[8], tmp8042[7], tmp8042[6], tmp8042[5], tmp8042[4], tmp8042[3], tmp8042[2], tmp8042[1], tmp8042[0]};
    assign tmp5464 = {tmp5463, const_461_0};
    assign tmp5481 = tmp5464 - tmp2887;
    assign tmp5482 = {tmp5481[16]};
    assign tmp5483 = {tmp5464[15]};
    assign tmp5484 = ~tmp5483;
    assign tmp5485 = tmp5482 ^ tmp5484;
    assign tmp5488 = tmp5485 ^ tmp6605;
    assign tmp5489 = tmp6100 & tmp5488;
    assign tmp5495 = {tmp3773[16]};
    assign tmp5506 = tmp2887 - tmp5464;
    assign tmp5507 = {tmp5506[16]};
    assign tmp5508 = {tmp2887[15]};
    assign tmp5510 = tmp5507 ^ tmp6605;
    assign tmp5513 = tmp5510 ^ tmp5484;
    assign tmp5514 = tmp2887 == tmp5464;
    assign tmp5515 = tmp5513 | tmp5514;
    assign tmp5516 = tmp3780 & tmp5515;
    assign tmp5517 = tmp5489 ? const_466_32767 : tmp5464;
    assign tmp5518 = tmp5516 ? _ver_out_tmp_62 : tmp5517;
    assign tmp5521 = tmp8058 - tmp5518;
    assign tmp5522 = {tmp5521[16]};
    assign tmp5525 = tmp5522 ^ tmp5173;
    assign tmp5526 = {tmp5518[15]};
    assign tmp5527 = ~tmp5526;
    assign tmp5528 = tmp5525 ^ tmp5527;
    assign tmp5550 = ~tmp5187;
    assign tmp5573 = {tmp5182[16]};
    assign tmp5576 = tmp5573 ^ tmp6605;
    assign tmp5580 = tmp2887 == tmp3253;
    assign tmp5581 = tmp5189 | tmp5580;
    assign tmp5587 = tmp8042 - tmp3307;
    assign tmp5588 = {tmp5587[16]};
    assign tmp5591 = tmp5588 ^ tmp3553;
    assign tmp5592 = {tmp3307[15]};
    assign tmp5593 = ~tmp5592;
    assign tmp5594 = tmp5591 ^ tmp5593;
    assign tmp5595 = tmp5528 & tmp5594;
    assign tmp5596 = {tmp8046[14], tmp8046[13], tmp8046[12], tmp8046[11], tmp8046[10], tmp8046[9], tmp8046[8], tmp8046[7], tmp8046[6], tmp8046[5], tmp8046[4], tmp8046[3], tmp8046[2], tmp8046[1], tmp8046[0]};
    assign tmp5597 = {tmp5596, const_475_0};
    assign tmp5603 = {tmp3867[16]};
    assign tmp5606 = tmp5603 ^ tmp6605;
    assign tmp5607 = {tmp8046[15]};
    assign tmp5609 = tmp5606 ^ tmp4623;
    assign tmp5614 = tmp5597 - tmp2887;
    assign tmp5615 = {tmp5614[16]};
    assign tmp5616 = {tmp5597[15]};
    assign tmp5617 = ~tmp5616;
    assign tmp5618 = tmp5615 ^ tmp5617;
    assign tmp5621 = tmp5618 ^ tmp6605;
    assign tmp5622 = tmp5609 & tmp5621;
    assign tmp5627 = tmp8046 - tmp2887;
    assign tmp5628 = {tmp5627[16]};
    assign tmp5631 = tmp5628 ^ tmp4623;
    assign tmp5634 = tmp5631 ^ tmp6605;
    assign tmp5639 = tmp2887 - tmp5597;
    assign tmp5640 = {tmp5639[16]};
    assign tmp5643 = tmp5640 ^ tmp6605;
    assign tmp5646 = tmp5643 ^ tmp5617;
    assign tmp5647 = tmp2887 == tmp5597;
    assign tmp5648 = tmp5646 | tmp5647;
    assign tmp5649 = tmp5634 & tmp5648;
    assign tmp5650 = tmp5622 ? const_480_32767 : tmp5597;
    assign tmp5651 = tmp5649 ? _ver_out_tmp_25 : tmp5650;
    assign tmp5654 = tmp8062 - tmp5651;
    assign tmp5655 = {tmp5654[16]};
    assign tmp5658 = tmp5655 ^ tmp3360;
    assign tmp5659 = {tmp5651[15]};
    assign tmp5660 = ~tmp5659;
    assign tmp5661 = tmp5658 ^ tmp5660;
    assign tmp5662 = tmp5595 & tmp5661;
    assign tmp5663 = {tmp8062[14], tmp8062[13], tmp8062[12], tmp8062[11], tmp8062[10], tmp8062[9], tmp8062[8], tmp8062[7], tmp8062[6], tmp8062[5], tmp8062[4], tmp8062[3], tmp8062[2], tmp8062[1], tmp8062[0]};
    assign tmp5669 = tmp2887 - tmp8062;
    assign tmp5670 = {tmp5669[16]};
    assign tmp5673 = tmp5670 ^ tmp6605;
    assign tmp5681 = tmp3327 - tmp2887;
    assign tmp5683 = {tmp3327[15]};
    assign tmp5689 = tmp4575 & tmp3351;
    assign tmp5694 = tmp8062 - tmp2887;
    assign tmp5701 = tmp3361 ^ tmp6605;
    assign tmp5706 = tmp2887 - tmp3327;
    assign tmp5707 = {tmp5706[16]};
    assign tmp5718 = tmp3379 ? _ver_out_tmp_66 : tmp5274;
    assign tmp5721 = tmp8046 - tmp5718;
    assign tmp5722 = {tmp5721[16]};
    assign tmp5725 = tmp5722 ^ tmp4623;
    assign tmp5726 = {tmp5718[15]};
    assign tmp5727 = ~tmp5726;
    assign tmp5728 = tmp5725 ^ tmp5727;
    assign tmp5729 = tmp5662 & tmp5728;
    assign tmp5730 = {tmp8050[14], tmp8050[13], tmp8050[12], tmp8050[11], tmp8050[10], tmp8050[9], tmp8050[8], tmp8050[7], tmp8050[6], tmp8050[5], tmp8050[4], tmp8050[3], tmp8050[2], tmp8050[1], tmp8050[0]};
    assign tmp5731 = {tmp5730, const_489_0};
    assign tmp5740 = tmp6390 ^ tmp6605;
    assign tmp5748 = tmp5731 - tmp2887;
    assign tmp5749 = {tmp5748[16]};
    assign tmp5752 = tmp5749 ^ tmp5779;
    assign tmp5755 = tmp5752 ^ tmp6605;
    assign tmp5756 = tmp4008 & tmp5755;
    assign tmp5768 = tmp4045 ^ tmp6605;
    assign tmp5773 = tmp2887 - tmp5731;
    assign tmp5774 = {tmp5773[16]};
    assign tmp5777 = tmp5774 ^ tmp6605;
    assign tmp5778 = {tmp5731[15]};
    assign tmp5779 = ~tmp5778;
    assign tmp5780 = tmp5777 ^ tmp5779;
    assign tmp5781 = tmp2887 == tmp5731;
    assign tmp5782 = tmp5780 | tmp5781;
    assign tmp5783 = tmp5768 & tmp5782;
    assign tmp5784 = tmp5756 ? const_494_32767 : tmp5731;
    assign tmp5785 = tmp5783 ? _ver_out_tmp_68 : tmp5784;
    assign tmp5788 = tmp8066 - tmp5785;
    assign tmp5789 = {tmp5788[16]};
    assign tmp5792 = tmp5789 ^ tmp4652;
    assign tmp5793 = {tmp5785[15]};
    assign tmp5794 = ~tmp5793;
    assign tmp5795 = tmp5792 ^ tmp5794;
    assign tmp5796 = tmp5729 & tmp5795;
    assign tmp5798 = {tmp5301, const_496_0};
    assign tmp5803 = tmp2887 - tmp8066;
    assign tmp5804 = {tmp5803[16]};
    assign tmp5815 = tmp5798 - tmp2887;
    assign tmp5817 = {tmp5798[15]};
    assign tmp5828 = tmp8066 - tmp2887;
    assign tmp5829 = {tmp5828[16]};
    assign tmp5835 = tmp3435 ^ tmp6605;
    assign tmp5840 = tmp2887 - tmp5798;
    assign tmp5844 = tmp5345 ^ tmp6605;
    assign tmp5846 = ~tmp5817;
    assign tmp5847 = tmp5844 ^ tmp5846;
    assign tmp5851 = tmp5327 ? const_501_32767 : tmp5798;
    assign tmp5855 = tmp8050 - tmp5356;
    assign tmp5856 = {tmp5855[16]};
    assign tmp5859 = tmp5856 ^ tmp4257;
    assign tmp5860 = {tmp5356[15]};
    assign tmp5861 = ~tmp5860;
    assign tmp5862 = tmp5859 ^ tmp5861;
    assign tmp5863 = tmp5796 & tmp5862;
    assign tmp5864 = {tmp8054[14], tmp8054[13], tmp8054[12], tmp8054[11], tmp8054[10], tmp8054[9], tmp8054[8], tmp8054[7], tmp8054[6], tmp8054[5], tmp8054[4], tmp8054[3], tmp8054[2], tmp8054[1], tmp8054[0]};
    assign tmp5865 = {tmp5864, const_503_0};
    assign tmp5871 = {tmp4135[16]};
    assign tmp5874 = tmp5871 ^ tmp6605;
    assign tmp5882 = tmp5865 - tmp2887;
    assign tmp5883 = {tmp5882[16]};
    assign tmp5886 = tmp5883 ^ tmp5913;
    assign tmp5889 = tmp5886 ^ tmp6605;
    assign tmp5890 = tmp4142 & tmp5889;
    assign tmp5899 = tmp6578 ^ tmp6543;
    assign tmp5907 = tmp2887 - tmp5865;
    assign tmp5908 = {tmp5907[16]};
    assign tmp5911 = tmp5908 ^ tmp6605;
    assign tmp5912 = {tmp5865[15]};
    assign tmp5913 = ~tmp5912;
    assign tmp5914 = tmp5911 ^ tmp5913;
    assign tmp5915 = tmp2887 == tmp5865;
    assign tmp5916 = tmp5914 | tmp5915;
    assign tmp5917 = tmp4182 & tmp5916;
    assign tmp5918 = tmp5890 ? const_508_32767 : tmp5865;
    assign tmp5919 = tmp5917 ? _ver_out_tmp_72 : tmp5918;
    assign tmp5922 = tmp8070 - tmp5919;
    assign tmp5923 = {tmp5922[16]};
    assign tmp5926 = tmp5923 ^ tmp3486;
    assign tmp5927 = {tmp5919[15]};
    assign tmp5928 = ~tmp5927;
    assign tmp5929 = tmp5926 ^ tmp5928;
    assign tmp5930 = tmp5863 & tmp5929;
    assign tmp5931 = {tmp8070[14], tmp8070[13], tmp8070[12], tmp8070[11], tmp8070[10], tmp8070[9], tmp8070[8], tmp8070[7], tmp8070[6], tmp8070[5], tmp8070[4], tmp8070[3], tmp8070[2], tmp8070[1], tmp8070[0]};
    assign tmp5932 = {tmp5931, const_510_0};
    assign tmp5941 = tmp4725 ^ tmp6605;
    assign tmp5952 = ~tmp5402;
    assign tmp5956 = tmp3496 ^ tmp6605;
    assign tmp5957 = tmp5395 & tmp5956;
    assign tmp5962 = tmp8070 - tmp2887;
    assign tmp5982 = tmp2887 == tmp5932;
    assign tmp5986 = tmp5435 ? _ver_out_tmp_74 : tmp3528;
    assign tmp5989 = tmp8054 - tmp5986;
    assign tmp5990 = {tmp5989[16]};
    assign tmp5993 = tmp5990 ^ tmp6543;
    assign tmp5994 = {tmp5986[15]};
    assign tmp5995 = ~tmp5994;
    assign tmp5996 = tmp5993 ^ tmp5995;
    assign tmp5997 = tmp5930 & tmp5996;
    assign tmp6072 = tmp6367 & tmp5997;
    assign tmp6083 = {tmp3719[16]};
    assign tmp6100 = tmp3737 ^ tmp3553;
    assign tmp6107 = {tmp6440[16]};
    assign tmp6109 = tmp3746 ^ tmp4016;
    assign tmp6127 = tmp3765 | tmp3766;
    assign tmp6128 = tmp3753 & tmp6127;
    assign tmp6149 = tmp3786 ^ tmp3788;
    assign tmp6152 = tmp6149 ^ tmp4016;
    assign tmp6159 = {tmp3798[16]};
    assign tmp6164 = ~tmp3760;
    assign tmp6165 = tmp3802 ^ tmp6164;
    assign tmp6167 = tmp6165 | tmp3766;
    assign tmp6168 = tmp3793 & tmp6167;
    assign tmp6169 = tmp6128 ? const_530_32767 : tmp3728;
    assign tmp6183 = tmp7435 & tmp8037;
    assign tmp6221 = _ver_out_tmp_81 == tmp8062;
    assign tmp6227 = tmp6221 ? tmp6864 : tmp5669;
    assign tmp6229 = {tmp5607, tmp5607};
    assign tmp6233 = {tmp3921, tmp6227};
    assign tmp6236 = {tmp3861[15], tmp3861[14], tmp3861[13], tmp3861[12], tmp3861[11], tmp3861[10], tmp3861[9], tmp3861[8], tmp3861[7], tmp3861[6], tmp3861[5], tmp3861[4], tmp3861[3], tmp3861[2], tmp3861[1], tmp3861[0]};
    assign tmp6253 = tmp6440 - tmp6227;
    assign tmp6257 = tmp3880 ^ tmp4016;
    assign tmp6260 = tmp6257 ^ tmp3922;
    assign tmp6261 = tmp5609 & tmp6260;
    assign tmp6270 = tmp3893 ^ tmp6312;
    assign tmp6273 = tmp6270 ^ tmp6605;
    assign tmp6276 = tmp6261 & tmp3901;
    assign tmp6294 = {tmp3919[17]};
    assign tmp6297 = tmp6294 ^ tmp3922;
    assign tmp6301 = tmp5634 & tmp3926;
    assign tmp6306 = tmp2887 - tmp6236;
    assign tmp6307 = {tmp6306[16]};
    assign tmp6310 = tmp6307 ^ tmp6605;
    assign tmp6312 = ~tmp3937;
    assign tmp6316 = tmp6301 & tmp3941;
    assign tmp6366 = ~tmp4784;
    assign tmp6367 = tmp5011 & tmp6366;
    assign tmp6369 = _ver_out_tmp_85 == tmp8066;
    assign tmp6377 = {tmp3988, tmp3988};
    assign tmp6381 = {tmp3991, tmp3987};
    assign tmp6382 = tmp3990 + tmp6381;
    assign tmp6390 = {tmp4001[16]};
    assign tmp6408 = tmp4017 ^ tmp4056;
    assign tmp6430 = {tmp4041[16]};
    assign tmp6440 = {tmp3742, const_554_0};
    assign tmp6462 = tmp2887 == tmp3996;
    assign tmp6463 = tmp4073 | tmp6462;
    assign tmp6517 = _ver_out_tmp_91 == tmp8070;
    assign tmp6523 = tmp6517 ? tmp6864 : tmp3480;
    assign tmp6526 = {tmp4123, tmp8054};
    assign tmp6542 = {tmp8054[15]};
    assign tmp6543 = ~tmp6542;
    assign tmp6549 = tmp6440 - tmp6523;
    assign tmp6550 = {tmp6549[17]};
    assign tmp6553 = tmp6550 ^ tmp4016;
    assign tmp6556 = tmp6553 ^ tmp4153;
    assign tmp6562 = tmp4130 - tmp2887;
    assign tmp6563 = {tmp6562[16]};
    assign tmp6566 = tmp6563 ^ tmp6608;
    assign tmp6569 = tmp6566 ^ tmp6605;
    assign tmp6577 = tmp8054 - tmp2887;
    assign tmp6578 = {tmp6577[16]};
    assign tmp6590 = {tmp4187[17]};
    assign tmp6591 = {tmp6523[16]};
    assign tmp6593 = tmp6590 ^ tmp4153;
    assign tmp6596 = tmp6593 ^ tmp4016;
    assign tmp6597 = tmp4182 & tmp6596;
    assign tmp6602 = tmp2887 - tmp4130;
    assign tmp6603 = {tmp6602[16]};
    assign tmp6605 = ~tmp5508;
    assign tmp6606 = tmp6603 ^ tmp6605;
    assign tmp6607 = {tmp4130[15]};
    assign tmp6608 = ~tmp6607;
    assign tmp6613 = tmp4170 ? const_569_32767 : tmp4130;
    assign tmp6633 = tmp6656 & tmp6657;
    assign tmp6634 = ~tmp4273;
    assign tmp6656 = tmp5209 & tmp4469;
    assign tmp6657 = ~tmp3658;
    assign tmp6665 = tmp6367 & tmp6690;
    assign tmp6690 = ~tmp5997;
    assign tmp6758 = {const_581_0, tmp11};
    assign tmp6759 = tmp586 ? tmp6758 : tmp2106;
    assign tmp6765 = {tmp2458[16]};
    assign tmp6772 = tmp15 == _ver_out_tmp_4;
    assign tmp6781 = tmp7154 ? tmp7163 : tmp2549;
    assign tmp6784 = tmp6759 - tmp6781;
    assign tmp6785 = {tmp6784[17]};
    assign tmp6786 = {tmp6759[16]};
    assign tmp6787 = ~tmp6786;
    assign tmp6788 = tmp6785 ^ tmp6787;
    assign tmp6791 = tmp6788 ^ tmp7173;
    assign tmp6808 = {const_594_0, const_594_0};
    assign tmp6813 = tmp2247 ? tmp7198 : tmp2492;
    assign tmp6825 = tmp376 ^ tmp6605;
    assign tmp6834 = {const_602_0, tmp16};
    assign tmp6838 = tmp6813 - tmp7225;
    assign tmp6839 = {tmp6838[17]};
    assign tmp6840 = {tmp6813[16]};
    assign tmp6841 = ~tmp6840;
    assign tmp6842 = tmp6839 ^ tmp6841;
    assign tmp6843 = {tmp7225[16]};
    assign tmp6844 = ~tmp6843;
    assign tmp6845 = tmp6842 ^ tmp6844;
    assign tmp6846 = tmp6791 & tmp6845;
    assign tmp6851 = tmp13 - tmp2887;
    assign tmp6864 = {tmp6808, const_607_32767};
    assign tmp6865 = tmp2885 ? tmp6864 : tmp7254;
    assign tmp6887 = tmp2581 ? tmp6864 : tmp7280;
    assign tmp6889 = {const_616_0, tmp17};
    assign tmp6890 = tmp2034 ? tmp6889 : tmp6887;
    assign tmp6893 = tmp7260 - tmp6890;
    assign tmp6894 = {tmp6893[17]};
    assign tmp6895 = {tmp7260[16]};
    assign tmp6896 = ~tmp6895;
    assign tmp6897 = tmp6894 ^ tmp6896;
    assign tmp6900 = tmp6897 ^ tmp7295;
    assign tmp6901 = tmp6846 & tmp6900;
    assign tmp6910 = tmp1790 ^ tmp2281;
    assign tmp6913 = tmp6910 ^ tmp6605;
    assign tmp6931 = ~tmp2041;
    assign tmp6935 = tmp2369 ^ tmp6605;
    assign tmp6936 = tmp18 == _ver_out_tmp_19;
    assign tmp6945 = tmp6935 ? tmp7346 : tmp2606;
    assign tmp6948 = tmp7321 - tmp6945;
    assign tmp6949 = {tmp6948[17]};
    assign tmp6950 = {tmp7321[16]};
    assign tmp6951 = ~tmp6950;
    assign tmp6952 = tmp6949 ^ tmp6951;
    assign tmp6953 = {tmp6945[16]};
    assign tmp6954 = ~tmp6953;
    assign tmp6955 = tmp6952 ^ tmp6954;
    assign tmp6956 = tmp6901 & tmp6955;
    assign tmp7020 = tmp7558 & tmp6956;
    assign tmp7031 = ~tmp2764;
    assign tmp7139 = {tmp6759[16], tmp6759[15], tmp6759[14], tmp6759[13], tmp6759[12], tmp6759[11], tmp6759[10], tmp6759[9], tmp6759[8], tmp6759[7], tmp6759[6], tmp6759[5], tmp6759[4], tmp6759[3], tmp6759[2], tmp6759[1]};
    assign tmp7140 = {tmp7139[15]};
    assign tmp7142 = {tmp7140, tmp7139};
    assign tmp7154 = tmp2807 ^ tmp6605;
    assign tmp7163 = {const_646_0, tmp15};
    assign tmp7167 = tmp6781 - tmp7142;
    assign tmp7168 = {tmp7167[17]};
    assign tmp7169 = {tmp7142[16]};
    assign tmp7170 = ~tmp7169;
    assign tmp7171 = tmp7168 ^ tmp7170;
    assign tmp7172 = {tmp6781[16]};
    assign tmp7173 = ~tmp7172;
    assign tmp7174 = tmp7171 ^ tmp7173;
    assign tmp7175 = tmp7142 == tmp6781;
    assign tmp7176 = tmp7174 | tmp7175;
    assign tmp7177 = tmp19 & tmp7176;
    assign tmp7185 = ~tmp1629;
    assign tmp7186 = tmp1665 ^ tmp7185;
    assign tmp7198 = {const_653_0, tmp12};
    assign tmp7200 = {tmp6813[16], tmp6813[15], tmp6813[14], tmp6813[13], tmp6813[12], tmp6813[11], tmp6813[10], tmp6813[9], tmp6813[8], tmp6813[7], tmp6813[6], tmp6813[5], tmp6813[4], tmp6813[3], tmp6813[2], tmp6813[1]};
    assign tmp7201 = {tmp7200[15]};
    assign tmp7203 = {tmp7201, tmp7200};
    assign tmp7225 = tmp6825 ? tmp6834 : tmp1092;
    assign tmp7228 = tmp7225 - tmp7203;
    assign tmp7229 = {tmp7228[17]};
    assign tmp7230 = {tmp7203[16]};
    assign tmp7231 = ~tmp7230;
    assign tmp7232 = tmp7229 ^ tmp7231;
    assign tmp7235 = tmp7232 ^ tmp6844;
    assign tmp7236 = tmp7203 == tmp7225;
    assign tmp7237 = tmp7235 | tmp7236;
    assign tmp7238 = tmp7177 & tmp7237;
    assign tmp7250 = tmp595 ^ tmp6605;
    assign tmp7254 = tmp2887 - tmp13;
    assign tmp7259 = {const_667_0, tmp13};
    assign tmp7260 = tmp7250 ? tmp7259 : tmp6865;
    assign tmp7261 = {tmp7260[16], tmp7260[15], tmp7260[14], tmp7260[13], tmp7260[12], tmp7260[11], tmp7260[10], tmp7260[9], tmp7260[8], tmp7260[7], tmp7260[6], tmp7260[5], tmp7260[4], tmp7260[3], tmp7260[2], tmp7260[1]};
    assign tmp7262 = {tmp7261[15]};
    assign tmp7264 = {tmp7262, tmp7261};
    assign tmp7280 = tmp2887 - tmp17;
    assign tmp7289 = tmp6890 - tmp7264;
    assign tmp7290 = {tmp7289[17]};
    assign tmp7291 = {tmp7264[16]};
    assign tmp7292 = ~tmp7291;
    assign tmp7293 = tmp7290 ^ tmp7292;
    assign tmp7294 = {tmp6890[16]};
    assign tmp7295 = ~tmp7294;
    assign tmp7296 = tmp7293 ^ tmp7295;
    assign tmp7297 = tmp7264 == tmp6890;
    assign tmp7298 = tmp7296 | tmp7297;
    assign tmp7299 = tmp7238 & tmp7298;
    assign tmp7320 = {const_681_0, tmp14};
    assign tmp7321 = tmp6913 ? tmp7320 : tmp2530;
    assign tmp7322 = {tmp7321[16], tmp7321[15], tmp7321[14], tmp7321[13], tmp7321[12], tmp7321[11], tmp7321[10], tmp7321[9], tmp7321[8], tmp7321[7], tmp7321[6], tmp7321[5], tmp7321[4], tmp7321[3], tmp7321[2], tmp7321[1]};
    assign tmp7323 = {tmp7322[15]};
    assign tmp7325 = {tmp7323, tmp7322};
    assign tmp7346 = {const_688_0, tmp18};
    assign tmp7350 = tmp6945 - tmp7325;
    assign tmp7351 = {tmp7350[17]};
    assign tmp7352 = {tmp7325[16]};
    assign tmp7353 = ~tmp7352;
    assign tmp7354 = tmp7351 ^ tmp7353;
    assign tmp7357 = tmp7354 ^ tmp6954;
    assign tmp7358 = tmp7325 == tmp6945;
    assign tmp7359 = tmp7357 | tmp7358;
    assign tmp7360 = tmp7299 & tmp7359;
    assign tmp7397 = {tmp11[15], tmp11[14], tmp11[13], tmp11[12], tmp11[11], tmp11[10], tmp11[9], tmp11[8], tmp11[7], tmp11[6], tmp11[5], tmp11[4], tmp11[3], tmp11[2], tmp11[1]};
    assign tmp7398 = {tmp7397[14]};
    assign tmp7400 = {tmp7398, tmp7397};
    assign tmp7419 = tmp7790 & tmp8038;
    assign tmp7420 = {tmp12[15], tmp12[14], tmp12[13], tmp12[12], tmp12[11], tmp12[10], tmp12[9], tmp12[8], tmp12[7], tmp12[6], tmp12[5], tmp12[4], tmp12[3], tmp12[2], tmp12[1]};
    assign tmp7421 = {tmp7420[14]};
    assign tmp7423 = {tmp7421, tmp7420};
    assign tmp7435 = tmp2681 & tmp7031;
    assign tmp7443 = {tmp13[15], tmp13[14], tmp13[13], tmp13[12], tmp13[11], tmp13[10], tmp13[9], tmp13[8], tmp13[7], tmp13[6], tmp13[5], tmp13[4], tmp13[3], tmp13[2], tmp13[1]};
    assign tmp7444 = {tmp7443[14]};
    assign tmp7446 = {tmp7444, tmp7443};
    assign tmp7466 = {tmp14[15], tmp14[14], tmp14[13], tmp14[12], tmp14[11], tmp14[10], tmp14[9], tmp14[8], tmp14[7], tmp14[6], tmp14[5], tmp14[4], tmp14[3], tmp14[2], tmp14[1]};
    assign tmp7467 = {tmp7466[14]};
    assign tmp7469 = {tmp7467, tmp7466};
    assign tmp7495 = tmp2887 - tmp15;
    assign tmp7511 = tmp293 ^ tmp7538;
    assign tmp7515 = tmp1340 & tmp1352;
    assign tmp7538 = ~tmp1347;
    assign tmp7558 = tmp7435 & tmp7785;
    assign tmp7564 = tmp7790 & tmp3196;
    assign tmp7565 = {tmp16[14], tmp16[13], tmp16[12], tmp16[11], tmp16[10], tmp16[9], tmp16[8], tmp16[7], tmp16[6], tmp16[5], tmp16[4], tmp16[3], tmp16[2], tmp16[1], tmp16[0]};
    assign tmp7572 = {tmp2565[16]};
    assign tmp7577 = ~tmp889;
    assign tmp7587 = tmp360 ^ tmp362;
    assign tmp7590 = tmp7587 ^ tmp6605;
    assign tmp7591 = tmp354 & tmp7590;
    assign tmp7596 = tmp16 - tmp2887;
    assign tmp7615 = tmp388 ^ tmp362;
    assign tmp7617 = tmp7615 | tmp392;
    assign tmp7618 = tmp6825 & tmp7617;
    assign tmp7620 = tmp7618 ? _ver_out_tmp_73 : tmp395;
    assign tmp7628 = ~tmp1113;
    assign tmp7641 = {tmp17[14], tmp17[13], tmp17[12], tmp17[11], tmp17[10], tmp17[9], tmp17[8], tmp17[7], tmp17[6], tmp17[5], tmp17[4], tmp17[3], tmp17[2], tmp17[1], tmp17[0]};
    assign tmp7651 = tmp1403 ^ tmp6605;
    assign tmp7654 = tmp7651 ^ tmp7675;
    assign tmp7660 = {tmp1414[16]};
    assign tmp7666 = tmp1418 ^ tmp6605;
    assign tmp7675 = ~tmp1429;
    assign tmp7684 = tmp2887 - tmp1397;
    assign tmp7688 = tmp1440 ^ tmp6605;
    assign tmp7692 = tmp2887 == tmp1397;
    assign tmp7695 = tmp1422 ? const_710_32767 : tmp1397;
    assign tmp7717 = {tmp18[14], tmp18[13], tmp18[12], tmp18[11], tmp18[10], tmp18[9], tmp18[8], tmp18[7], tmp18[6], tmp18[5], tmp18[4], tmp18[3], tmp18[2], tmp18[1], tmp18[0]};
    assign tmp7718 = {tmp7717, const_712_0};
    assign tmp7735 = tmp7718 - tmp2887;
    assign tmp7736 = {tmp7735[16]};
    assign tmp7738 = ~tmp7765;
    assign tmp7739 = tmp7736 ^ tmp7738;
    assign tmp7742 = tmp7739 ^ tmp6605;
    assign tmp7743 = tmp2006 & tmp7742;
    assign tmp7760 = tmp2887 - tmp7718;
    assign tmp7761 = {tmp7760[16]};
    assign tmp7764 = tmp7761 ^ tmp6605;
    assign tmp7765 = {tmp7718[15]};
    assign tmp7767 = tmp7764 ^ tmp7738;
    assign tmp7768 = tmp2887 == tmp7718;
    assign tmp7769 = tmp7767 | tmp7768;
    assign tmp7770 = tmp6935 & tmp7769;
    assign tmp7771 = tmp7743 ? const_717_32767 : tmp7718;
    assign tmp7772 = tmp7770 ? _ver_out_tmp_2 : tmp7771;
    assign tmp7785 = ~tmp8037;
    assign tmp7790 = tmp7809 & tmp7360;
    assign tmp7809 = tmp7558 & tmp7827;
    assign tmp7810 = ~tmp7360;
    assign tmp7818 = tmp4971 & tmp8130;
    assign tmp7827 = ~tmp6956;
    assign tmp7830 = tmp7809 & tmp7810;
    assign tmp7863 = tmp73 ? const_6_0 : tmp11;
    assign tmp7864 = tmp273 ? tmp195 : tmp7863;
    assign tmp7865 = tmp427 ? tmp13 : tmp7864;
    assign tmp7866 = tmp873 ? tmp616 : tmp7865;
    assign tmp7867 = tmp1110 ? tmp2474 : tmp7866;
    assign tmp7868 = tmp1464 ? tmp195 : tmp7867;
    assign tmp7869 = tmp1561 ? tmp12 : tmp7868;
    assign tmp7870 = tmp2081 ? tmp1689 : tmp7869;
    assign tmp7871 = tmp2126 ? tmp2474 : tmp7870;
    assign tmp7872 = tmp2826 ? tmp2474 : tmp7871;
    assign tmp7873 = tmp3145 ? tmp3602 : tmp7872;
    assign tmp7874 = tmp3215 ? tmp8042 : tmp7873;
    assign tmp7875 = tmp3694 ? tmp8058 : tmp7874;
    assign tmp7876 = tmp4413 ? tmp8058 : tmp7875;
    assign tmp7877 = tmp4886 ? tmp3602 : tmp7876;
    assign tmp7878 = tmp5219 ? tmp8042 : tmp7877;
    assign tmp7879 = tmp6072 ? tmp8058 : tmp7878;
    assign tmp7880 = tmp7020 ? tmp15 : tmp7879;
    assign tmp7881 = tmp7419 ? tmp7400 : tmp7880;
    assign tmp7882 = tmp73 ? const_7_2 : tmp12;
    assign tmp7883 = tmp273 ? tmp262 : tmp7882;
    assign tmp7884 = tmp427 ? tmp14 : tmp7883;
    assign tmp7885 = tmp873 ? tmp737 : tmp7884;
    assign tmp7886 = tmp1110 ? tmp2870 : tmp7885;
    assign tmp7887 = tmp1166 ? tmp11 : tmp7886;
    assign tmp7888 = tmp1561 ? tmp11 : tmp7887;
    assign tmp7889 = tmp2081 ? tmp11 : tmp7888;
    assign tmp7890 = tmp2826 ? tmp2870 : tmp7889;
    assign tmp7891 = tmp3145 ? tmp2948 : tmp7890;
    assign tmp7892 = tmp3215 ? tmp8046 : tmp7891;
    assign tmp7893 = tmp3694 ? tmp8062 : tmp7892;
    assign tmp7894 = tmp4413 ? tmp8062 : tmp7893;
    assign tmp7895 = tmp4886 ? tmp2948 : tmp7894;
    assign tmp7896 = tmp5219 ? tmp8046 : tmp7895;
    assign tmp7897 = tmp6072 ? tmp8062 : tmp7896;
    assign tmp7898 = tmp7020 ? tmp16 : tmp7897;
    assign tmp7899 = tmp7419 ? tmp7423 : tmp7898;
    assign tmp7900 = tmp73 ? const_8_1 : tmp13;
    assign tmp7901 = tmp119 ? tmp11 : tmp7900;
    assign tmp7902 = tmp427 ? tmp11 : tmp7901;
    assign tmp7903 = tmp873 ? tmp11 : tmp7902;
    assign tmp7904 = tmp1464 ? tmp1313 : tmp7903;
    assign tmp7905 = tmp1561 ? tmp14 : tmp7904;
    assign tmp7906 = tmp2081 ? tmp1814 : tmp7905;
    assign tmp7907 = tmp2126 ? tmp2512 : tmp7906;
    assign tmp7908 = tmp2826 ? tmp2512 : tmp7907;
    assign tmp7909 = tmp3145 ? tmp4890 : tmp7908;
    assign tmp7910 = tmp3215 ? tmp8050 : tmp7909;
    assign tmp7911 = tmp3694 ? tmp8066 : tmp7910;
    assign tmp7912 = tmp4413 ? tmp8066 : tmp7911;
    assign tmp7913 = tmp4886 ? tmp4890 : tmp7912;
    assign tmp7914 = tmp5219 ? tmp8050 : tmp7913;
    assign tmp7915 = tmp6072 ? tmp8066 : tmp7914;
    assign tmp7916 = tmp7020 ? tmp17 : tmp7915;
    assign tmp7917 = tmp7419 ? tmp7446 : tmp7916;
    assign tmp7918 = tmp73 ? const_9_0 : tmp14;
    assign tmp7919 = tmp119 ? tmp12 : tmp7918;
    assign tmp7920 = tmp427 ? tmp12 : tmp7919;
    assign tmp7921 = tmp873 ? tmp12 : tmp7920;
    assign tmp7922 = tmp1166 ? tmp13 : tmp7921;
    assign tmp7923 = tmp1561 ? tmp13 : tmp7922;
    assign tmp7924 = tmp2081 ? tmp13 : tmp7923;
    assign tmp7925 = tmp2826 ? tmp2531 : tmp7924;
    assign tmp7926 = tmp3145 ? tmp2982 : tmp7925;
    assign tmp7927 = tmp3215 ? tmp8054 : tmp7926;
    assign tmp7928 = tmp3694 ? tmp8070 : tmp7927;
    assign tmp7929 = tmp4413 ? tmp8070 : tmp7928;
    assign tmp7930 = tmp4886 ? tmp2982 : tmp7929;
    assign tmp7931 = tmp5219 ? tmp8054 : tmp7930;
    assign tmp7932 = tmp6072 ? tmp8070 : tmp7931;
    assign tmp7933 = tmp7020 ? tmp18 : tmp7932;
    assign tmp7934 = tmp7419 ? tmp7469 : tmp7933;
    assign tmp7935 = tmp73 ? const_10_0 : tmp15;
    assign tmp7936 = tmp273 ? tmp329 : tmp7935;
    assign tmp7937 = tmp427 ? tmp17 : tmp7936;
    assign tmp7938 = tmp873 ? tmp858 : tmp7937;
    assign tmp7939 = tmp1110 ? tmp2550 : tmp7938;
    assign tmp7940 = tmp1464 ? tmp329 : tmp7939;
    assign tmp7941 = tmp1561 ? tmp16 : tmp7940;
    assign tmp7942 = tmp2081 ? tmp1939 : tmp7941;
    assign tmp7943 = tmp2126 ? tmp2550 : tmp7942;
    assign tmp7944 = tmp3145 ? tmp8058 : tmp7943;
    assign tmp7945 = tmp3215 ? tmp3307 : tmp7944;
    assign tmp7946 = tmp3694 ? tmp3810 : tmp7945;
    assign tmp7947 = tmp4413 ? tmp8042 : tmp7946;
    assign tmp7948 = tmp4886 ? tmp8058 : tmp7947;
    assign tmp7949 = tmp5219 ? tmp3307 : tmp7948;
    assign tmp7950 = tmp6072 ? tmp3810 : tmp7949;
    assign tmp7951 = tmp7020 ? tmp11 : tmp7950;
    assign tmp7952 = tmp7564 ? tmp329 : tmp7951;
    assign tmp7953 = tmp73 ? const_11_0 : tmp16;
    assign tmp7954 = tmp273 ? tmp7620 : tmp7953;
    assign tmp7955 = tmp427 ? tmp18 : tmp7954;
    assign tmp7956 = tmp873 ? tmp979 : tmp7955;
    assign tmp7957 = tmp1110 ? tmp2569 : tmp7956;
    assign tmp7958 = tmp1166 ? tmp15 : tmp7957;
    assign tmp7959 = tmp1561 ? tmp15 : tmp7958;
    assign tmp7960 = tmp2081 ? tmp15 : tmp7959;
    assign tmp7961 = tmp3145 ? tmp8062 : tmp7960;
    assign tmp7962 = tmp3215 ? tmp5718 : tmp7961;
    assign tmp7963 = tmp3694 ? tmp3944 : tmp7962;
    assign tmp7964 = tmp4413 ? tmp8046 : tmp7963;
    assign tmp7965 = tmp4886 ? tmp8062 : tmp7964;
    assign tmp7966 = tmp5219 ? tmp5718 : tmp7965;
    assign tmp7967 = tmp6072 ? tmp3944 : tmp7966;
    assign tmp7968 = tmp7020 ? tmp12 : tmp7967;
    assign tmp7969 = tmp7564 ? tmp7620 : tmp7968;
    assign tmp7970 = tmp73 ? const_12_0 : tmp17;
    assign tmp7971 = tmp119 ? tmp15 : tmp7970;
    assign tmp7972 = tmp427 ? tmp15 : tmp7971;
    assign tmp7973 = tmp873 ? tmp15 : tmp7972;
    assign tmp7974 = tmp1464 ? tmp1451 : tmp7973;
    assign tmp7975 = tmp1561 ? tmp18 : tmp7974;
    assign tmp7976 = tmp2081 ? tmp2064 : tmp7975;
    assign tmp7977 = tmp2126 ? tmp2588 : tmp7976;
    assign tmp7978 = tmp3145 ? tmp8066 : tmp7977;
    assign tmp7979 = tmp3215 ? tmp5356 : tmp7978;
    assign tmp7980 = tmp3694 ? tmp4078 : tmp7979;
    assign tmp7981 = tmp4413 ? tmp8050 : tmp7980;
    assign tmp7982 = tmp4886 ? tmp8066 : tmp7981;
    assign tmp7983 = tmp5219 ? tmp5356 : tmp7982;
    assign tmp7984 = tmp6072 ? tmp4078 : tmp7983;
    assign tmp7985 = tmp7020 ? tmp13 : tmp7984;
    assign tmp7986 = tmp7564 ? tmp1451 : tmp7985;
    assign tmp7987 = tmp73 ? const_13_1 : tmp18;
    assign tmp7988 = tmp119 ? tmp16 : tmp7987;
    assign tmp7989 = tmp427 ? tmp16 : tmp7988;
    assign tmp7990 = tmp873 ? tmp16 : tmp7989;
    assign tmp7991 = tmp1166 ? tmp17 : tmp7990;
    assign tmp7992 = tmp1561 ? tmp17 : tmp7991;
    assign tmp7993 = tmp2081 ? tmp17 : tmp7992;
    assign tmp7994 = tmp3145 ? tmp8070 : tmp7993;
    assign tmp7995 = tmp3215 ? tmp5986 : tmp7994;
    assign tmp7996 = tmp3694 ? tmp4212 : tmp7995;
    assign tmp7997 = tmp4413 ? tmp8054 : tmp7996;
    assign tmp7998 = tmp4886 ? tmp8070 : tmp7997;
    assign tmp7999 = tmp5219 ? tmp5986 : tmp7998;
    assign tmp8000 = tmp6072 ? tmp4212 : tmp7999;
    assign tmp8001 = tmp7020 ? tmp14 : tmp8000;
    assign tmp8002 = tmp7564 ? tmp7772 : tmp8001;
    assign tmp8003 = tmp73 ? const_14_0 : tmp19;
    assign tmp8004 = tmp459 ? tmp19 : tmp8003;
    assign tmp8005 = tmp1141 ? tmp19 : tmp8004;
    assign tmp8006 = tmp2775 ? const_292_0 : tmp8005;
    assign tmp8007 = tmp2826 ? const_296_0 : tmp8006;
    assign tmp8008 = tmp3397 ? const_318_0 : tmp8007;
    assign tmp8009 = tmp3694 ? const_348_0 : tmp8008;
    assign tmp8010 = tmp4413 ? const_402_0 : tmp8009;
    assign tmp8011 = tmp5013 ? const_432_0 : tmp8010;
    assign tmp8012 = tmp6072 ? const_518_1 : tmp8011;
    assign tmp8013 = tmp6665 ? const_572_0 : tmp8012;
    assign tmp8014 = const_782_0 ? const_574_0 : tmp8013;
    assign tmp8015 = tmp7020 ? const_632_1 : tmp8014;
    assign tmp8016 = tmp7790 ? const_690_1 : tmp8015;
    assign tmp8017 = tmp7830 ? tmp19 : tmp8016;
    assign tmp8018 = const_783_0 ? tmp19 : tmp8017;
    assign tmp8019 = tmp459 ? const_17_0 : my_calculator_out_z;
    assign tmp8020 = tmp1141 ? const_118_0 : tmp8019;
    assign tmp8021 = tmp2775 ? const_291_15 : tmp8020;
    assign tmp8022 = tmp2826 ? const_295_8 : tmp8021;
    assign tmp8023 = tmp3397 ? const_317_1 : tmp8022;
    assign tmp8024 = tmp3694 ? const_347_4 : tmp8023;
    assign tmp8025 = tmp4413 ? const_401_6 : tmp8024;
    assign tmp8026 = tmp5013 ? const_431_2 : tmp8025;
    assign tmp8027 = tmp6072 ? const_517_5 : tmp8026;
    assign tmp8028 = tmp6665 ? const_571_0 : tmp8027;
    assign tmp8029 = const_784_0 ? const_573_0 : tmp8028;
    assign tmp8030 = tmp7020 ? const_631_6 : tmp8029;
    assign tmp8031 = tmp7790 ? const_689_3 : tmp8030;
    assign tmp8032 = tmp7830 ? const_719_0 : tmp8031;
    assign tmp8033 = const_781_0 ? const_720_0 : tmp8032;
    assign tmp8034 = tmp2681 ? tmp2287 : const_721_0;
    assign tmp8035 = tmp2681 ? tmp2374 : const_722_0;
    assign tmp8036 = tmp2681 ? tmp2399 : const_723_0;
    assign tmp8037 = tmp2681 ? tmp2412 : const_724_0;
    assign tmp8038 = tmp2681 ? tmp2430 : const_725_0;
    assign tmp8041 = tmp2561 ? tmp2474 : tmp2887;
    assign tmp8042 = tmp2736 ? tmp11 : tmp8041;
    assign tmp8045 = tmp2561 ? tmp2870 : tmp2887;
    assign tmp8046 = tmp2736 ? tmp12 : tmp8045;
    assign tmp8049 = tmp2561 ? tmp2512 : tmp2887;
    assign tmp8050 = tmp2736 ? tmp13 : tmp8049;
    assign tmp8053 = tmp2561 ? tmp2531 : tmp2887;
    assign tmp8054 = tmp2736 ? tmp14 : tmp8053;
    assign tmp8057 = tmp2561 ? tmp2550 : tmp2887;
    assign tmp8058 = tmp2736 ? tmp15 : tmp8057;
    assign tmp8061 = tmp2561 ? tmp2569 : tmp2887;
    assign tmp8062 = tmp2736 ? tmp16 : tmp8061;
    assign tmp8065 = tmp2561 ? tmp2588 : tmp2887;
    assign tmp8066 = tmp2736 ? tmp17 : tmp8065;
    assign tmp8069 = tmp2561 ? tmp2607 : tmp2887;
    assign tmp8070 = tmp2736 ? tmp18 : tmp8069;
    assign tmp8074 = tmp8071 == tmp1179;
    assign tmp8076 = {tmp6808, const_744_2};
    assign tmp8077 = tmp8071 == tmp8076;
    assign tmp8078 = tmp8074 | tmp8077;
    assign tmp8080 = {tmp6808, const_746_3};
    assign tmp8081 = tmp8071 == tmp8080;
    assign tmp8082 = tmp8078 | tmp8081;
    assign tmp8083 = tmp8071 == const_748_15;
    assign tmp8084 = tmp8082 | tmp8083;
    assign tmp8087 = tmp8071 == tmp520;
    assign tmp8090 = tmp8071 == tmp523;
    assign tmp8091 = tmp8087 | tmp8090;
    assign tmp8095 = tmp8091 | tmp8105;
    assign tmp8099 = tmp8095 | tmp8109;
    assign tmp8101 = tmp8099 | tmp8083;
    assign tmp8102 = tmp8071 == const_758_8;
    assign tmp8104 = {const_760_0, const_759_6};
    assign tmp8105 = tmp8071 == tmp8104;
    assign tmp8106 = tmp8102 | tmp8105;
    assign tmp8108 = {const_762_0, const_761_7};
    assign tmp8109 = tmp8071 == tmp8108;
    assign tmp8110 = tmp8106 | tmp8109;
    assign tmp8112 = tmp8110 | tmp8083;
    assign tmp8114 = tmp5 == tmp8;
    assign tmp8117 = {tmp6808, const_764_1};
    assign tmp8118 = my_calculator_ctrl == tmp8117;
    assign tmp8120 = tmp10 & tmp8118;
    assign tmp8126 = tmp8141 & tmp1113;
    assign tmp8129 = my_calculator_ctrl == tmp2209;
    assign tmp8130 = ~tmp8118;
    assign tmp8138 = tmp8141 & tmp7628;
    assign tmp8141 = tmp10 & tmp8130;
    assign tmp8144 = tmp8138 & tmp8129;
    assign tmp8149 = ~tmp8129;
    assign tmp8156 = tmp8138 & tmp8149;
    assign tmp8157 = tmp8120 ? const_766_2 : my_calculator_ctrl;
    assign tmp8158 = tmp8126 ? const_770_3 : tmp8157;
    assign tmp8159 = tmp8144 ? const_773_1 : tmp8158;
    assign tmp8160 = tmp8156 ? const_775_1 : tmp8159;
    assign tmp8161 = tmp8120 ? const_767_15 : my_calculator_in_y;
    assign tmp8162 = tmp8144 ? const_774_15 : my_calculator_in_x;
    assign tmp8163 = tmp8156 ? const_776_15 : tmp8162;
    assign tmp8164 = tmp8144 ? my_calculator_out_z : tmp8071;

    // Registers
    always @(posedge clk)
    begin
        begin
            my_calculator_ctrl <= tmp8160;
            my_calculator_in_x <= tmp8163;
            my_calculator_in_y <= tmp8161;
            my_calculator_out_z <= tmp8033;
            tmp0 <= tmp4;
            tmp5 <= tmp8;
            tmp7 <= tmp10;
            tmp11 <= tmp7881;
            tmp12 <= tmp7899;
            tmp13 <= tmp7917;
            tmp14 <= tmp7934;
            tmp15 <= tmp7952;
            tmp16 <= tmp7969;
            tmp17 <= tmp7986;
            tmp18 <= tmp8002;
            tmp19 <= tmp8018;
            tmp8071 <= tmp8164;
        end
    end

endmodule

